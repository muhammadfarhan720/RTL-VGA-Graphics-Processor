
module pika_name_g(
	input clock,
	input [9:0] address,
	output reg [7:0] data_out
);

reg [7:0] mem [0:1023];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 8'b00001111;
	mem[1] = 8'b00001111;
	mem[2] = 8'b00001110;
	mem[3] = 8'b00001101;
	mem[4] = 8'b00001111;
	mem[5] = 8'b00001111;
	mem[6] = 8'b00001111;
	mem[7] = 8'b00001111;
	mem[8] = 8'b00001111;
	mem[9] = 8'b00001111;
	mem[10] = 8'b00001111;
	mem[11] = 8'b00001111;
	mem[12] = 8'b00001111;
	mem[13] = 8'b00001111;
	mem[14] = 8'b00001111;
	mem[15] = 8'b00001111;
	mem[16] = 8'b00001111;
	mem[17] = 8'b00001111;
	mem[18] = 8'b00001111;
	mem[19] = 8'b00001111;
	mem[20] = 8'b00001111;
	mem[21] = 8'b00001111;
	mem[22] = 8'b00001111;
	mem[23] = 8'b00001111;
	mem[24] = 8'b00001111;
	mem[25] = 8'b00001111;
	mem[26] = 8'b00001111;
	mem[27] = 8'b00001111;
	mem[28] = 8'b00001111;
	mem[29] = 8'b00001111;
	mem[30] = 8'b00001111;
	mem[31] = 8'b00001111;
	mem[32] = 8'b00001111;
	mem[33] = 8'b00001111;
	mem[34] = 8'b00001111;
	mem[35] = 8'b00001111;
	mem[36] = 8'b00001111;
	mem[37] = 8'b00001111;
	mem[38] = 8'b00001111;
	mem[39] = 8'b00001111;
	mem[40] = 8'b00001111;
	mem[41] = 8'b00001111;
	mem[42] = 8'b00001111;
	mem[43] = 8'b00001111;
	mem[44] = 8'b00001111;
	mem[45] = 8'b00001111;
	mem[46] = 8'b00001111;
	mem[47] = 8'b00001111;
	mem[48] = 8'b00001111;
	mem[49] = 8'b00001111;
	mem[50] = 8'b00001111;
	mem[51] = 8'b00001111;
	mem[52] = 8'b00001111;
	mem[53] = 8'b00001111;
	mem[54] = 8'b00001111;
	mem[55] = 8'b00001111;
	mem[56] = 8'b00001111;
	mem[57] = 8'b00001111;
	mem[58] = 8'b00001111;
	mem[59] = 8'b00001111;
	mem[60] = 8'b00001111;
	mem[61] = 8'b00001111;
	mem[62] = 8'b00001110;
	mem[63] = 8'b00001011;
	mem[64] = 8'b00001111;
	mem[65] = 8'b00001111;
	mem[66] = 8'b00001010;
	mem[67] = 8'b00001100;
	mem[68] = 8'b00001011;
	mem[69] = 8'b00001010;
	mem[70] = 8'b00001010;
	mem[71] = 8'b00001100;
	mem[72] = 8'b00001111;
	mem[73] = 8'b00001111;
	mem[74] = 8'b00001111;
	mem[75] = 8'b00001111;
	mem[76] = 8'b00001111;
	mem[77] = 8'b00001111;
	mem[78] = 8'b00001111;
	mem[79] = 8'b00001111;
	mem[80] = 8'b00001111;
	mem[81] = 8'b00001111;
	mem[82] = 8'b00001111;
	mem[83] = 8'b00001111;
	mem[84] = 8'b00001111;
	mem[85] = 8'b00001111;
	mem[86] = 8'b00001111;
	mem[87] = 8'b00001111;
	mem[88] = 8'b00001111;
	mem[89] = 8'b00001111;
	mem[90] = 8'b00001111;
	mem[91] = 8'b00001111;
	mem[92] = 8'b00001111;
	mem[93] = 8'b00001111;
	mem[94] = 8'b00001111;
	mem[95] = 8'b00001111;
	mem[96] = 8'b00001111;
	mem[97] = 8'b00001111;
	mem[98] = 8'b00001111;
	mem[99] = 8'b00001111;
	mem[100] = 8'b00001111;
	mem[101] = 8'b00001111;
	mem[102] = 8'b00001111;
	mem[103] = 8'b00001111;
	mem[104] = 8'b00001111;
	mem[105] = 8'b00001111;
	mem[106] = 8'b00001111;
	mem[107] = 8'b00001111;
	mem[108] = 8'b00001111;
	mem[109] = 8'b00001111;
	mem[110] = 8'b00001111;
	mem[111] = 8'b00001111;
	mem[112] = 8'b00001111;
	mem[113] = 8'b00001111;
	mem[114] = 8'b00001111;
	mem[115] = 8'b00001111;
	mem[116] = 8'b00001111;
	mem[117] = 8'b00001111;
	mem[118] = 8'b00001111;
	mem[119] = 8'b00001100;
	mem[120] = 8'b00001010;
	mem[121] = 8'b00001010;
	mem[122] = 8'b00001111;
	mem[123] = 8'b00001111;
	mem[124] = 8'b00001111;
	mem[125] = 8'b00001010;
	mem[126] = 8'b00001100;
	mem[127] = 8'b00001001;
	mem[128] = 8'b00001111;
	mem[129] = 8'b00001111;
	mem[130] = 8'b00001010;
	mem[131] = 8'b00001100;
	mem[132] = 8'b00001100;
	mem[133] = 8'b00001100;
	mem[134] = 8'b00001100;
	mem[135] = 8'b00001100;
	mem[136] = 8'b00001010;
	mem[137] = 8'b00001111;
	mem[138] = 8'b00001111;
	mem[139] = 8'b00001101;
	mem[140] = 8'b00001010;
	mem[141] = 8'b00001010;
	mem[142] = 8'b00001100;
	mem[143] = 8'b00001111;
	mem[144] = 8'b00001111;
	mem[145] = 8'b00001011;
	mem[146] = 8'b00001100;
	mem[147] = 8'b00001110;
	mem[148] = 8'b00001111;
	mem[149] = 8'b00001111;
	mem[150] = 8'b00001101;
	mem[151] = 8'b00001010;
	mem[152] = 8'b00001111;
	mem[153] = 8'b00001111;
	mem[154] = 8'b00001111;
	mem[155] = 8'b00001111;
	mem[156] = 8'b00001111;
	mem[157] = 8'b00001111;
	mem[158] = 8'b00001111;
	mem[159] = 8'b00001110;
	mem[160] = 8'b00001111;
	mem[161] = 8'b00001110;
	mem[162] = 8'b00001111;
	mem[163] = 8'b00001111;
	mem[164] = 8'b00001111;
	mem[165] = 8'b00001111;
	mem[166] = 8'b00001111;
	mem[167] = 8'b00001111;
	mem[168] = 8'b00001111;
	mem[169] = 8'b00001111;
	mem[170] = 8'b00001111;
	mem[171] = 8'b00001111;
	mem[172] = 8'b00001111;
	mem[173] = 8'b00001110;
	mem[174] = 8'b00001011;
	mem[175] = 8'b00001011;
	mem[176] = 8'b00001111;
	mem[177] = 8'b00001111;
	mem[178] = 8'b00001111;
	mem[179] = 8'b00001010;
	mem[180] = 8'b00001011;
	mem[181] = 8'b00001001;
	mem[182] = 8'b00001111;
	mem[183] = 8'b00001010;
	mem[184] = 8'b00001100;
	mem[185] = 8'b00001001;
	mem[186] = 8'b00001111;
	mem[187] = 8'b00001111;
	mem[188] = 8'b00001111;
	mem[189] = 8'b00001011;
	mem[190] = 8'b00001100;
	mem[191] = 8'b00001001;
	mem[192] = 8'b00001111;
	mem[193] = 8'b00001101;
	mem[194] = 8'b00001100;
	mem[195] = 8'b00001100;
	mem[196] = 8'b00001000;
	mem[197] = 8'b00001001;
	mem[198] = 8'b00001001;
	mem[199] = 8'b00001100;
	mem[200] = 8'b00001010;
	mem[201] = 8'b00001111;
	mem[202] = 8'b00001111;
	mem[203] = 8'b00001010;
	mem[204] = 8'b00001100;
	mem[205] = 8'b00001011;
	mem[206] = 8'b00001101;
	mem[207] = 8'b00001111;
	mem[208] = 8'b00001100;
	mem[209] = 8'b00001100;
	mem[210] = 8'b00001100;
	mem[211] = 8'b00001011;
	mem[212] = 8'b00001111;
	mem[213] = 8'b00001010;
	mem[214] = 8'b00001100;
	mem[215] = 8'b00001100;
	mem[216] = 8'b00001001;
	mem[217] = 8'b00001111;
	mem[218] = 8'b00001111;
	mem[219] = 8'b00001111;
	mem[220] = 8'b00001111;
	mem[221] = 8'b00001111;
	mem[222] = 8'b00001100;
	mem[223] = 8'b00001011;
	mem[224] = 8'b00001011;
	mem[225] = 8'b00001001;
	mem[226] = 8'b00001111;
	mem[227] = 8'b00001111;
	mem[228] = 8'b00001111;
	mem[229] = 8'b00001111;
	mem[230] = 8'b00001100;
	mem[231] = 8'b00001010;
	mem[232] = 8'b00001011;
	mem[233] = 8'b00001100;
	mem[234] = 8'b00001001;
	mem[235] = 8'b00001111;
	mem[236] = 8'b00001111;
	mem[237] = 8'b00001010;
	mem[238] = 8'b00001100;
	mem[239] = 8'b00001010;
	mem[240] = 8'b00001111;
	mem[241] = 8'b00001111;
	mem[242] = 8'b00001111;
	mem[243] = 8'b00001100;
	mem[244] = 8'b00001100;
	mem[245] = 8'b00001001;
	mem[246] = 8'b00001111;
	mem[247] = 8'b00001100;
	mem[248] = 8'b00001100;
	mem[249] = 8'b00001001;
	mem[250] = 8'b00001111;
	mem[251] = 8'b00001111;
	mem[252] = 8'b00001101;
	mem[253] = 8'b00001100;
	mem[254] = 8'b00001100;
	mem[255] = 8'b00001011;
	mem[256] = 8'b00001111;
	mem[257] = 8'b00001010;
	mem[258] = 8'b00001100;
	mem[259] = 8'b00001100;
	mem[260] = 8'b00001010;
	mem[261] = 8'b00001101;
	mem[262] = 8'b00001010;
	mem[263] = 8'b00001100;
	mem[264] = 8'b00001010;
	mem[265] = 8'b00001111;
	mem[266] = 8'b00001111;
	mem[267] = 8'b00001010;
	mem[268] = 8'b00001100;
	mem[269] = 8'b00001001;
	mem[270] = 8'b00001111;
	mem[271] = 8'b00001111;
	mem[272] = 8'b00001010;
	mem[273] = 8'b00001100;
	mem[274] = 8'b00001001;
	mem[275] = 8'b00001011;
	mem[276] = 8'b00001011;
	mem[277] = 8'b00001100;
	mem[278] = 8'b00001100;
	mem[279] = 8'b00001001;
	mem[280] = 8'b00001101;
	mem[281] = 8'b00001111;
	mem[282] = 8'b00001111;
	mem[283] = 8'b00001111;
	mem[284] = 8'b00001111;
	mem[285] = 8'b00001100;
	mem[286] = 8'b00001100;
	mem[287] = 8'b00001100;
	mem[288] = 8'b00001100;
	mem[289] = 8'b00001011;
	mem[290] = 8'b00001111;
	mem[291] = 8'b00001111;
	mem[292] = 8'b00001110;
	mem[293] = 8'b00001010;
	mem[294] = 8'b00001100;
	mem[295] = 8'b00001100;
	mem[296] = 8'b00001010;
	mem[297] = 8'b00001010;
	mem[298] = 8'b00001000;
	mem[299] = 8'b00001111;
	mem[300] = 8'b00001111;
	mem[301] = 8'b00001011;
	mem[302] = 8'b00001100;
	mem[303] = 8'b00001001;
	mem[304] = 8'b00001111;
	mem[305] = 8'b00001111;
	mem[306] = 8'b00001011;
	mem[307] = 8'b00001100;
	mem[308] = 8'b00001100;
	mem[309] = 8'b00001100;
	mem[310] = 8'b00001011;
	mem[311] = 8'b00001100;
	mem[312] = 8'b00001011;
	mem[313] = 8'b00001110;
	mem[314] = 8'b00001111;
	mem[315] = 8'b00001111;
	mem[316] = 8'b00001010;
	mem[317] = 8'b00001100;
	mem[318] = 8'b00001010;
	mem[319] = 8'b00001111;
	mem[320] = 8'b00001111;
	mem[321] = 8'b00001010;
	mem[322] = 8'b00001100;
	mem[323] = 8'b00001100;
	mem[324] = 8'b00001100;
	mem[325] = 8'b00001100;
	mem[326] = 8'b00001100;
	mem[327] = 8'b00001100;
	mem[328] = 8'b00001000;
	mem[329] = 8'b00001111;
	mem[330] = 8'b00001101;
	mem[331] = 8'b00001100;
	mem[332] = 8'b00001100;
	mem[333] = 8'b00001001;
	mem[334] = 8'b00001111;
	mem[335] = 8'b00001111;
	mem[336] = 8'b00001011;
	mem[337] = 8'b00001100;
	mem[338] = 8'b00001011;
	mem[339] = 8'b00001100;
	mem[340] = 8'b00001100;
	mem[341] = 8'b00001010;
	mem[342] = 8'b00001010;
	mem[343] = 8'b00001111;
	mem[344] = 8'b00001111;
	mem[345] = 8'b00001111;
	mem[346] = 8'b00001111;
	mem[347] = 8'b00001111;
	mem[348] = 8'b00001101;
	mem[349] = 8'b00001011;
	mem[350] = 8'b00001100;
	mem[351] = 8'b00001001;
	mem[352] = 8'b00001100;
	mem[353] = 8'b00001100;
	mem[354] = 8'b00001100;
	mem[355] = 8'b00001110;
	mem[356] = 8'b00001011;
	mem[357] = 8'b00001100;
	mem[358] = 8'b00001010;
	mem[359] = 8'b00001010;
	mem[360] = 8'b00001111;
	mem[361] = 8'b00001111;
	mem[362] = 8'b00001111;
	mem[363] = 8'b00001111;
	mem[364] = 8'b00001100;
	mem[365] = 8'b00001100;
	mem[366] = 8'b00001100;
	mem[367] = 8'b00001001;
	mem[368] = 8'b00001010;
	mem[369] = 8'b00001010;
	mem[370] = 8'b00001011;
	mem[371] = 8'b00001100;
	mem[372] = 8'b00001001;
	mem[373] = 8'b00001111;
	mem[374] = 8'b00001010;
	mem[375] = 8'b00001100;
	mem[376] = 8'b00001001;
	mem[377] = 8'b00001111;
	mem[378] = 8'b00001111;
	mem[379] = 8'b00001111;
	mem[380] = 8'b00001010;
	mem[381] = 8'b00001100;
	mem[382] = 8'b00001001;
	mem[383] = 8'b00001111;
	mem[384] = 8'b00001110;
	mem[385] = 8'b00001100;
	mem[386] = 8'b00001100;
	mem[387] = 8'b00001001;
	mem[388] = 8'b00001001;
	mem[389] = 8'b00001010;
	mem[390] = 8'b00001001;
	mem[391] = 8'b00001001;
	mem[392] = 8'b00001111;
	mem[393] = 8'b00001111;
	mem[394] = 8'b00001010;
	mem[395] = 8'b00001100;
	mem[396] = 8'b00001010;
	mem[397] = 8'b00001110;
	mem[398] = 8'b00001111;
	mem[399] = 8'b00001011;
	mem[400] = 8'b00001100;
	mem[401] = 8'b00001100;
	mem[402] = 8'b00001100;
	mem[403] = 8'b00001011;
	mem[404] = 8'b00001001;
	mem[405] = 8'b00001111;
	mem[406] = 8'b00001111;
	mem[407] = 8'b00001111;
	mem[408] = 8'b00001111;
	mem[409] = 8'b00001111;
	mem[410] = 8'b00001111;
	mem[411] = 8'b00001101;
	mem[412] = 8'b00001011;
	mem[413] = 8'b00001100;
	mem[414] = 8'b00001010;
	mem[415] = 8'b00001101;
	mem[416] = 8'b00001011;
	mem[417] = 8'b00001100;
	mem[418] = 8'b00001001;
	mem[419] = 8'b00001010;
	mem[420] = 8'b00001100;
	mem[421] = 8'b00001010;
	mem[422] = 8'b00001101;
	mem[423] = 8'b00001111;
	mem[424] = 8'b00001111;
	mem[425] = 8'b00001111;
	mem[426] = 8'b00001111;
	mem[427] = 8'b00001111;
	mem[428] = 8'b00001010;
	mem[429] = 8'b00001100;
	mem[430] = 8'b00001100;
	mem[431] = 8'b00001100;
	mem[432] = 8'b00001100;
	mem[433] = 8'b00001101;
	mem[434] = 8'b00001100;
	mem[435] = 8'b00001100;
	mem[436] = 8'b00001001;
	mem[437] = 8'b00001111;
	mem[438] = 8'b00001011;
	mem[439] = 8'b00001100;
	mem[440] = 8'b00001001;
	mem[441] = 8'b00001111;
	mem[442] = 8'b00001111;
	mem[443] = 8'b00001101;
	mem[444] = 8'b00001100;
	mem[445] = 8'b00001100;
	mem[446] = 8'b00001001;
	mem[447] = 8'b00001111;
	mem[448] = 8'b00001011;
	mem[449] = 8'b00001100;
	mem[450] = 8'b00001011;
	mem[451] = 8'b00001100;
	mem[452] = 8'b00001111;
	mem[453] = 8'b00001111;
	mem[454] = 8'b00001111;
	mem[455] = 8'b00001111;
	mem[456] = 8'b00001111;
	mem[457] = 8'b00001111;
	mem[458] = 8'b00001011;
	mem[459] = 8'b00001100;
	mem[460] = 8'b00001001;
	mem[461] = 8'b00001111;
	mem[462] = 8'b00001111;
	mem[463] = 8'b00001010;
	mem[464] = 8'b00001100;
	mem[465] = 8'b00001100;
	mem[466] = 8'b00001100;
	mem[467] = 8'b00001010;
	mem[468] = 8'b00001110;
	mem[469] = 8'b00001111;
	mem[470] = 8'b00001111;
	mem[471] = 8'b00001111;
	mem[472] = 8'b00001111;
	mem[473] = 8'b00001111;
	mem[474] = 8'b00001101;
	mem[475] = 8'b00001011;
	mem[476] = 8'b00001100;
	mem[477] = 8'b00001100;
	mem[478] = 8'b00001010;
	mem[479] = 8'b00001010;
	mem[480] = 8'b00001100;
	mem[481] = 8'b00001100;
	mem[482] = 8'b00001001;
	mem[483] = 8'b00001010;
	mem[484] = 8'b00001100;
	mem[485] = 8'b00001001;
	mem[486] = 8'b00001111;
	mem[487] = 8'b00001111;
	mem[488] = 8'b00001111;
	mem[489] = 8'b00001110;
	mem[490] = 8'b00001111;
	mem[491] = 8'b00001111;
	mem[492] = 8'b00001011;
	mem[493] = 8'b00001100;
	mem[494] = 8'b00001001;
	mem[495] = 8'b00001010;
	mem[496] = 8'b00001010;
	mem[497] = 8'b00001001;
	mem[498] = 8'b00001100;
	mem[499] = 8'b00001011;
	mem[500] = 8'b00001100;
	mem[501] = 8'b00001101;
	mem[502] = 8'b00001100;
	mem[503] = 8'b00001100;
	mem[504] = 8'b00001011;
	mem[505] = 8'b00001111;
	mem[506] = 8'b00001110;
	mem[507] = 8'b00001010;
	mem[508] = 8'b00001100;
	mem[509] = 8'b00001010;
	mem[510] = 8'b00001110;
	mem[511] = 8'b00001111;
	mem[512] = 8'b00001010;
	mem[513] = 8'b00001100;
	mem[514] = 8'b00001001;
	mem[515] = 8'b00001111;
	mem[516] = 8'b00001111;
	mem[517] = 8'b00001111;
	mem[518] = 8'b00001111;
	mem[519] = 8'b00001111;
	mem[520] = 8'b00001111;
	mem[521] = 8'b00001100;
	mem[522] = 8'b00001100;
	mem[523] = 8'b00001100;
	mem[524] = 8'b00001010;
	mem[525] = 8'b00001111;
	mem[526] = 8'b00001110;
	mem[527] = 8'b00001100;
	mem[528] = 8'b00001100;
	mem[529] = 8'b00001000;
	mem[530] = 8'b00001010;
	mem[531] = 8'b00001100;
	mem[532] = 8'b00001010;
	mem[533] = 8'b00001101;
	mem[534] = 8'b00001111;
	mem[535] = 8'b00001111;
	mem[536] = 8'b00001111;
	mem[537] = 8'b00001101;
	mem[538] = 8'b00001011;
	mem[539] = 8'b00001100;
	mem[540] = 8'b00001011;
	mem[541] = 8'b00001010;
	mem[542] = 8'b00001010;
	mem[543] = 8'b00001010;
	mem[544] = 8'b00001011;
	mem[545] = 8'b00001100;
	mem[546] = 8'b00001001;
	mem[547] = 8'b00001010;
	mem[548] = 8'b00001100;
	mem[549] = 8'b00001011;
	mem[550] = 8'b00001010;
	mem[551] = 8'b00001010;
	mem[552] = 8'b00001010;
	mem[553] = 8'b00001011;
	mem[554] = 8'b00001011;
	mem[555] = 8'b00001011;
	mem[556] = 8'b00001100;
	mem[557] = 8'b00001011;
	mem[558] = 8'b00001101;
	mem[559] = 8'b00001111;
	mem[560] = 8'b00001111;
	mem[561] = 8'b00001010;
	mem[562] = 8'b00001100;
	mem[563] = 8'b00001001;
	mem[564] = 8'b00001111;
	mem[565] = 8'b00001110;
	mem[566] = 8'b00001100;
	mem[567] = 8'b00001100;
	mem[568] = 8'b00001010;
	mem[569] = 8'b00001010;
	mem[570] = 8'b00001011;
	mem[571] = 8'b00001100;
	mem[572] = 8'b00001011;
	mem[573] = 8'b00001010;
	mem[574] = 8'b00001111;
	mem[575] = 8'b00001111;
	mem[576] = 8'b00001001;
	mem[577] = 8'b00001010;
	mem[578] = 8'b00001001;
	mem[579] = 8'b00001111;
	mem[580] = 8'b00001111;
	mem[581] = 8'b00001111;
	mem[582] = 8'b00001111;
	mem[583] = 8'b00001111;
	mem[584] = 8'b00001111;
	mem[585] = 8'b00001001;
	mem[586] = 8'b00001100;
	mem[587] = 8'b00001010;
	mem[588] = 8'b00001111;
	mem[589] = 8'b00001111;
	mem[590] = 8'b00001010;
	mem[591] = 8'b00001100;
	mem[592] = 8'b00001010;
	mem[593] = 8'b00001111;
	mem[594] = 8'b00001101;
	mem[595] = 8'b00001010;
	mem[596] = 8'b00001100;
	mem[597] = 8'b00001011;
	mem[598] = 8'b00001100;
	mem[599] = 8'b00001111;
	mem[600] = 8'b00001111;
	mem[601] = 8'b00001010;
	mem[602] = 8'b00001100;
	mem[603] = 8'b00001001;
	mem[604] = 8'b00001101;
	mem[605] = 8'b00001111;
	mem[606] = 8'b00001111;
	mem[607] = 8'b00001111;
	mem[608] = 8'b00001010;
	mem[609] = 8'b00001100;
	mem[610] = 8'b00001010;
	mem[611] = 8'b00001101;
	mem[612] = 8'b00001001;
	mem[613] = 8'b00001100;
	mem[614] = 8'b00001100;
	mem[615] = 8'b00001100;
	mem[616] = 8'b00001011;
	mem[617] = 8'b00001001;
	mem[618] = 8'b00001010;
	mem[619] = 8'b00001010;
	mem[620] = 8'b00001100;
	mem[621] = 8'b00001001;
	mem[622] = 8'b00001111;
	mem[623] = 8'b00001111;
	mem[624] = 8'b00001101;
	mem[625] = 8'b00001100;
	mem[626] = 8'b00001100;
	mem[627] = 8'b00001001;
	mem[628] = 8'b00001111;
	mem[629] = 8'b00001111;
	mem[630] = 8'b00001010;
	mem[631] = 8'b00001011;
	mem[632] = 8'b00001100;
	mem[633] = 8'b00001100;
	mem[634] = 8'b00001100;
	mem[635] = 8'b00001010;
	mem[636] = 8'b00001010;
	mem[637] = 8'b00001111;
	mem[638] = 8'b00001111;
	mem[639] = 8'b00001111;
	mem[640] = 8'b00001111;
	mem[641] = 8'b00001111;
	mem[642] = 8'b00001111;
	mem[643] = 8'b00001111;
	mem[644] = 8'b00001111;
	mem[645] = 8'b00001111;
	mem[646] = 8'b00001111;
	mem[647] = 8'b00001111;
	mem[648] = 8'b00001111;
	mem[649] = 8'b00001111;
	mem[650] = 8'b00001010;
	mem[651] = 8'b00001010;
	mem[652] = 8'b00001111;
	mem[653] = 8'b00001111;
	mem[654] = 8'b00001100;
	mem[655] = 8'b00001001;
	mem[656] = 8'b00001001;
	mem[657] = 8'b00001111;
	mem[658] = 8'b00001111;
	mem[659] = 8'b00001110;
	mem[660] = 8'b00001001;
	mem[661] = 8'b00001001;
	mem[662] = 8'b00001110;
	mem[663] = 8'b00001111;
	mem[664] = 8'b00001111;
	mem[665] = 8'b00001110;
	mem[666] = 8'b00001001;
	mem[667] = 8'b00001101;
	mem[668] = 8'b00001111;
	mem[669] = 8'b00001111;
	mem[670] = 8'b00001111;
	mem[671] = 8'b00001111;
	mem[672] = 8'b00001101;
	mem[673] = 8'b00001010;
	mem[674] = 8'b00001011;
	mem[675] = 8'b00001111;
	mem[676] = 8'b00001111;
	mem[677] = 8'b00001101;
	mem[678] = 8'b00001011;
	mem[679] = 8'b00001011;
	mem[680] = 8'b00001110;
	mem[681] = 8'b00001111;
	mem[682] = 8'b00001111;
	mem[683] = 8'b00001011;
	mem[684] = 8'b00001001;
	mem[685] = 8'b00001011;
	mem[686] = 8'b00001111;
	mem[687] = 8'b00001111;
	mem[688] = 8'b00001111;
	mem[689] = 8'b00001011;
	mem[690] = 8'b00001001;
	mem[691] = 8'b00001110;
	mem[692] = 8'b00001111;
	mem[693] = 8'b00001111;
	mem[694] = 8'b00001111;
	mem[695] = 8'b00001101;
	mem[696] = 8'b00001010;
	mem[697] = 8'b00001010;
	mem[698] = 8'b00001010;
	mem[699] = 8'b00001111;
	mem[700] = 8'b00001111;
	mem[701] = 8'b00001111;
	mem[702] = 8'b00001111;
	mem[703] = 8'b00001111;
	mem[704] = 8'b00000000;
	mem[705] = 8'b00000000;
	mem[706] = 8'b00000000;
	mem[707] = 8'b00000000;
	mem[708] = 8'b00000000;
	mem[709] = 8'b00000000;
	mem[710] = 8'b00000000;
	mem[711] = 8'b00000000;
	mem[712] = 8'b00000000;
	mem[713] = 8'b00000000;
	mem[714] = 8'b00000000;
	mem[715] = 8'b00000000;
	mem[716] = 8'b00000000;
	mem[717] = 8'b00000000;
	mem[718] = 8'b00000000;
	mem[719] = 8'b00000000;
	mem[720] = 8'b00000000;
	mem[721] = 8'b00000000;
	mem[722] = 8'b00000000;
	mem[723] = 8'b00000000;
	mem[724] = 8'b00000000;
	mem[725] = 8'b00000000;
	mem[726] = 8'b00000000;
	mem[727] = 8'b00000000;
	mem[728] = 8'b00000000;
	mem[729] = 8'b00000000;
	mem[730] = 8'b00000000;
	mem[731] = 8'b00000000;
	mem[732] = 8'b00000000;
	mem[733] = 8'b00000000;
	mem[734] = 8'b00000000;
	mem[735] = 8'b00000000;
	mem[736] = 8'b00000000;
	mem[737] = 8'b00000000;
	mem[738] = 8'b00000000;
	mem[739] = 8'b00000000;
	mem[740] = 8'b00000000;
	mem[741] = 8'b00000000;
	mem[742] = 8'b00000000;
	mem[743] = 8'b00000000;
	mem[744] = 8'b00000000;
	mem[745] = 8'b00000000;
	mem[746] = 8'b00000000;
	mem[747] = 8'b00000000;
	mem[748] = 8'b00000000;
	mem[749] = 8'b00000000;
	mem[750] = 8'b00000000;
	mem[751] = 8'b00000000;
	mem[752] = 8'b00000000;
	mem[753] = 8'b00000000;
	mem[754] = 8'b00000000;
	mem[755] = 8'b00000000;
	mem[756] = 8'b00000000;
	mem[757] = 8'b00000000;
	mem[758] = 8'b00000000;
	mem[759] = 8'b00000000;
	mem[760] = 8'b00000000;
	mem[761] = 8'b00000000;
	mem[762] = 8'b00000000;
	mem[763] = 8'b00000000;
	mem[764] = 8'b00000000;
	mem[765] = 8'b00000000;
	mem[766] = 8'b00000000;
	mem[767] = 8'b00000000;
	mem[768] = 8'b00000000;
	mem[769] = 8'b00000000;
	mem[770] = 8'b00000000;
	mem[771] = 8'b00000000;
	mem[772] = 8'b00000000;
	mem[773] = 8'b00000000;
	mem[774] = 8'b00000000;
	mem[775] = 8'b00000000;
	mem[776] = 8'b00000000;
	mem[777] = 8'b00000000;
	mem[778] = 8'b00000000;
	mem[779] = 8'b00000000;
	mem[780] = 8'b00000000;
	mem[781] = 8'b00000000;
	mem[782] = 8'b00000000;
	mem[783] = 8'b00000000;
	mem[784] = 8'b00000000;
	mem[785] = 8'b00000000;
	mem[786] = 8'b00000000;
	mem[787] = 8'b00000000;
	mem[788] = 8'b00000000;
	mem[789] = 8'b00000000;
	mem[790] = 8'b00000000;
	mem[791] = 8'b00000000;
	mem[792] = 8'b00000000;
	mem[793] = 8'b00000000;
	mem[794] = 8'b00000000;
	mem[795] = 8'b00000000;
	mem[796] = 8'b00000000;
	mem[797] = 8'b00000000;
	mem[798] = 8'b00000000;
	mem[799] = 8'b00000000;
	mem[800] = 8'b00000000;
	mem[801] = 8'b00000000;
	mem[802] = 8'b00000000;
	mem[803] = 8'b00000000;
	mem[804] = 8'b00000000;
	mem[805] = 8'b00000000;
	mem[806] = 8'b00000000;
	mem[807] = 8'b00000000;
	mem[808] = 8'b00000000;
	mem[809] = 8'b00000000;
	mem[810] = 8'b00000000;
	mem[811] = 8'b00000000;
	mem[812] = 8'b00000000;
	mem[813] = 8'b00000000;
	mem[814] = 8'b00000000;
	mem[815] = 8'b00000000;
	mem[816] = 8'b00000000;
	mem[817] = 8'b00000000;
	mem[818] = 8'b00000000;
	mem[819] = 8'b00000000;
	mem[820] = 8'b00000000;
	mem[821] = 8'b00000000;
	mem[822] = 8'b00000000;
	mem[823] = 8'b00000000;
	mem[824] = 8'b00000000;
	mem[825] = 8'b00000000;
	mem[826] = 8'b00000000;
	mem[827] = 8'b00000000;
	mem[828] = 8'b00000000;
	mem[829] = 8'b00000000;
	mem[830] = 8'b00000000;
	mem[831] = 8'b00000000;
	mem[832] = 8'b00000000;
	mem[833] = 8'b00000000;
	mem[834] = 8'b00000000;
	mem[835] = 8'b00000000;
	mem[836] = 8'b00000000;
	mem[837] = 8'b00000000;
	mem[838] = 8'b00000000;
	mem[839] = 8'b00000000;
	mem[840] = 8'b00000000;
	mem[841] = 8'b00000000;
	mem[842] = 8'b00000000;
	mem[843] = 8'b00000000;
	mem[844] = 8'b00000000;
	mem[845] = 8'b00000000;
	mem[846] = 8'b00000000;
	mem[847] = 8'b00000000;
	mem[848] = 8'b00000000;
	mem[849] = 8'b00000000;
	mem[850] = 8'b00000000;
	mem[851] = 8'b00000000;
	mem[852] = 8'b00000000;
	mem[853] = 8'b00000000;
	mem[854] = 8'b00000000;
	mem[855] = 8'b00000000;
	mem[856] = 8'b00000000;
	mem[857] = 8'b00000000;
	mem[858] = 8'b00000000;
	mem[859] = 8'b00000000;
	mem[860] = 8'b00000000;
	mem[861] = 8'b00000000;
	mem[862] = 8'b00000000;
	mem[863] = 8'b00000000;
	mem[864] = 8'b00000000;
	mem[865] = 8'b00000000;
	mem[866] = 8'b00000000;
	mem[867] = 8'b00000000;
	mem[868] = 8'b00000000;
	mem[869] = 8'b00000000;
	mem[870] = 8'b00000000;
	mem[871] = 8'b00000000;
	mem[872] = 8'b00000000;
	mem[873] = 8'b00000000;
	mem[874] = 8'b00000000;
	mem[875] = 8'b00000000;
	mem[876] = 8'b00000000;
	mem[877] = 8'b00000000;
	mem[878] = 8'b00000000;
	mem[879] = 8'b00000000;
	mem[880] = 8'b00000000;
	mem[881] = 8'b00000000;
	mem[882] = 8'b00000000;
	mem[883] = 8'b00000000;
	mem[884] = 8'b00000000;
	mem[885] = 8'b00000000;
	mem[886] = 8'b00000000;
	mem[887] = 8'b00000000;
	mem[888] = 8'b00000000;
	mem[889] = 8'b00000000;
	mem[890] = 8'b00000000;
	mem[891] = 8'b00000000;
	mem[892] = 8'b00000000;
	mem[893] = 8'b00000000;
	mem[894] = 8'b00000000;
	mem[895] = 8'b00000000;
	mem[896] = 8'b00000000;
	mem[897] = 8'b00000000;
	mem[898] = 8'b00000000;
	mem[899] = 8'b00000000;
	mem[900] = 8'b00000000;
	mem[901] = 8'b00000000;
	mem[902] = 8'b00000000;
	mem[903] = 8'b00000000;
	mem[904] = 8'b00000000;
	mem[905] = 8'b00000000;
	mem[906] = 8'b00000000;
	mem[907] = 8'b00000000;
	mem[908] = 8'b00000000;
	mem[909] = 8'b00000000;
	mem[910] = 8'b00000000;
	mem[911] = 8'b00000000;
	mem[912] = 8'b00000000;
	mem[913] = 8'b00000000;
	mem[914] = 8'b00000000;
	mem[915] = 8'b00000000;
	mem[916] = 8'b00000000;
	mem[917] = 8'b00000000;
	mem[918] = 8'b00000000;
	mem[919] = 8'b00000000;
	mem[920] = 8'b00000000;
	mem[921] = 8'b00000000;
	mem[922] = 8'b00000000;
	mem[923] = 8'b00000000;
	mem[924] = 8'b00000000;
	mem[925] = 8'b00000000;
	mem[926] = 8'b00000000;
	mem[927] = 8'b00000000;
	mem[928] = 8'b00000000;
	mem[929] = 8'b00000000;
	mem[930] = 8'b00000000;
	mem[931] = 8'b00000000;
	mem[932] = 8'b00000000;
	mem[933] = 8'b00000000;
	mem[934] = 8'b00000000;
	mem[935] = 8'b00000000;
	mem[936] = 8'b00000000;
	mem[937] = 8'b00000000;
	mem[938] = 8'b00000000;
	mem[939] = 8'b00000000;
	mem[940] = 8'b00000000;
	mem[941] = 8'b00000000;
	mem[942] = 8'b00000000;
	mem[943] = 8'b00000000;
	mem[944] = 8'b00000000;
	mem[945] = 8'b00000000;
	mem[946] = 8'b00000000;
	mem[947] = 8'b00000000;
	mem[948] = 8'b00000000;
	mem[949] = 8'b00000000;
	mem[950] = 8'b00000000;
	mem[951] = 8'b00000000;
	mem[952] = 8'b00000000;
	mem[953] = 8'b00000000;
	mem[954] = 8'b00000000;
	mem[955] = 8'b00000000;
	mem[956] = 8'b00000000;
	mem[957] = 8'b00000000;
	mem[958] = 8'b00000000;
	mem[959] = 8'b00000000;
	mem[960] = 8'b00000000;
	mem[961] = 8'b00000000;
	mem[962] = 8'b00000000;
	mem[963] = 8'b00000000;
	mem[964] = 8'b00000000;
	mem[965] = 8'b00000000;
	mem[966] = 8'b00000000;
	mem[967] = 8'b00000000;
	mem[968] = 8'b00000000;
	mem[969] = 8'b00000000;
	mem[970] = 8'b00000000;
	mem[971] = 8'b00000000;
	mem[972] = 8'b00000000;
	mem[973] = 8'b00000000;
	mem[974] = 8'b00000000;
	mem[975] = 8'b00000000;
	mem[976] = 8'b00000000;
	mem[977] = 8'b00000000;
	mem[978] = 8'b00000000;
	mem[979] = 8'b00000000;
	mem[980] = 8'b00000000;
	mem[981] = 8'b00000000;
	mem[982] = 8'b00000000;
	mem[983] = 8'b00000000;
	mem[984] = 8'b00000000;
	mem[985] = 8'b00000000;
	mem[986] = 8'b00000000;
	mem[987] = 8'b00000000;
	mem[988] = 8'b00000000;
	mem[989] = 8'b00000000;
	mem[990] = 8'b00000000;
	mem[991] = 8'b00000000;
	mem[992] = 8'b00000000;
	mem[993] = 8'b00000000;
	mem[994] = 8'b00000000;
	mem[995] = 8'b00000000;
	mem[996] = 8'b00000000;
	mem[997] = 8'b00000000;
	mem[998] = 8'b00000000;
	mem[999] = 8'b00000000;
	mem[1000] = 8'b00000000;
	mem[1001] = 8'b00000000;
	mem[1002] = 8'b00000000;
	mem[1003] = 8'b00000000;
	mem[1004] = 8'b00000000;
	mem[1005] = 8'b00000000;
	mem[1006] = 8'b00000000;
	mem[1007] = 8'b00000000;
	mem[1008] = 8'b00000000;
	mem[1009] = 8'b00000000;
	mem[1010] = 8'b00000000;
	mem[1011] = 8'b00000000;
	mem[1012] = 8'b00000000;
	mem[1013] = 8'b00000000;
	mem[1014] = 8'b00000000;
	mem[1015] = 8'b00000000;
	mem[1016] = 8'b00000000;
	mem[1017] = 8'b00000000;
	mem[1018] = 8'b00000000;
	mem[1019] = 8'b00000000;
	mem[1020] = 8'b00000000;
	mem[1021] = 8'b00000000;
	mem[1022] = 8'b00000000;
	mem[1023] = 8'b00000000;
end
endmodule
