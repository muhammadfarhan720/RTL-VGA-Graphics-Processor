
module attack_rom_g(
	input clock,
	input [10:0] address,
	output reg [7:0] data_out
);

reg [7:0] mem [0:2047];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 8'b00001111;
	mem[1] = 8'b00001111;
	mem[2] = 8'b00001111;
	mem[3] = 8'b00001111;
	mem[4] = 8'b00001111;
	mem[5] = 8'b00001111;
	mem[6] = 8'b00001111;
	mem[7] = 8'b00001111;
	mem[8] = 8'b00001111;
	mem[9] = 8'b00001111;
	mem[10] = 8'b00001111;
	mem[11] = 8'b00001111;
	mem[12] = 8'b00001111;
	mem[13] = 8'b00001111;
	mem[14] = 8'b00001111;
	mem[15] = 8'b00001111;
	mem[16] = 8'b00001100;
	mem[17] = 8'b00001011;
	mem[18] = 8'b00001011;
	mem[19] = 8'b00001011;
	mem[20] = 8'b00001011;
	mem[21] = 8'b00001011;
	mem[22] = 8'b00001011;
	mem[23] = 8'b00001011;
	mem[24] = 8'b00001100;
	mem[25] = 8'b00001111;
	mem[26] = 8'b00001111;
	mem[27] = 8'b00001111;
	mem[28] = 8'b00001111;
	mem[29] = 8'b00001111;
	mem[30] = 8'b00001111;
	mem[31] = 8'b00001111;
	mem[32] = 8'b00001111;
	mem[33] = 8'b00001111;
	mem[34] = 8'b00001111;
	mem[35] = 8'b00001111;
	mem[36] = 8'b00001111;
	mem[37] = 8'b00001111;
	mem[38] = 8'b00001111;
	mem[39] = 8'b00001111;
	mem[40] = 8'b00001111;
	mem[41] = 8'b00001111;
	mem[42] = 8'b00001111;
	mem[43] = 8'b00001111;
	mem[44] = 8'b00001111;
	mem[45] = 8'b00001111;
	mem[46] = 8'b00001111;
	mem[47] = 8'b00001111;
	mem[48] = 8'b00001111;
	mem[49] = 8'b00001111;
	mem[50] = 8'b00001111;
	mem[51] = 8'b00001111;
	mem[52] = 8'b00001111;
	mem[53] = 8'b00001111;
	mem[54] = 8'b00001111;
	mem[55] = 8'b00001111;
	mem[56] = 8'b00001111;
	mem[57] = 8'b00001111;
	mem[58] = 8'b00001111;
	mem[59] = 8'b00001111;
	mem[60] = 8'b00001111;
	mem[61] = 8'b00001111;
	mem[62] = 8'b00001111;
	mem[63] = 8'b00001111;
	mem[64] = 8'b00001111;
	mem[65] = 8'b00001111;
	mem[66] = 8'b00001111;
	mem[67] = 8'b00001111;
	mem[68] = 8'b00001111;
	mem[69] = 8'b00001111;
	mem[70] = 8'b00001111;
	mem[71] = 8'b00001111;
	mem[72] = 8'b00001111;
	mem[73] = 8'b00001111;
	mem[74] = 8'b00001111;
	mem[75] = 8'b00001111;
	mem[76] = 8'b00001111;
	mem[77] = 8'b00001111;
	mem[78] = 8'b00001011;
	mem[79] = 8'b00001010;
	mem[80] = 8'b00001011;
	mem[81] = 8'b00001011;
	mem[82] = 8'b00001011;
	mem[83] = 8'b00001011;
	mem[84] = 8'b00001011;
	mem[85] = 8'b00001011;
	mem[86] = 8'b00001011;
	mem[87] = 8'b00001011;
	mem[88] = 8'b00001011;
	mem[89] = 8'b00001010;
	mem[90] = 8'b00001100;
	mem[91] = 8'b00001111;
	mem[92] = 8'b00001111;
	mem[93] = 8'b00001111;
	mem[94] = 8'b00001111;
	mem[95] = 8'b00001111;
	mem[96] = 8'b00001111;
	mem[97] = 8'b00001111;
	mem[98] = 8'b00001111;
	mem[99] = 8'b00001111;
	mem[100] = 8'b00001111;
	mem[101] = 8'b00001111;
	mem[102] = 8'b00001111;
	mem[103] = 8'b00001111;
	mem[104] = 8'b00001111;
	mem[105] = 8'b00001111;
	mem[106] = 8'b00001111;
	mem[107] = 8'b00001111;
	mem[108] = 8'b00001111;
	mem[109] = 8'b00001111;
	mem[110] = 8'b00001111;
	mem[111] = 8'b00001111;
	mem[112] = 8'b00001111;
	mem[113] = 8'b00001111;
	mem[114] = 8'b00001111;
	mem[115] = 8'b00001111;
	mem[116] = 8'b00001111;
	mem[117] = 8'b00001111;
	mem[118] = 8'b00001111;
	mem[119] = 8'b00001111;
	mem[120] = 8'b00001111;
	mem[121] = 8'b00001111;
	mem[122] = 8'b00001111;
	mem[123] = 8'b00001111;
	mem[124] = 8'b00001111;
	mem[125] = 8'b00001111;
	mem[126] = 8'b00001111;
	mem[127] = 8'b00001111;
	mem[128] = 8'b00001111;
	mem[129] = 8'b00001111;
	mem[130] = 8'b00001111;
	mem[131] = 8'b00001111;
	mem[132] = 8'b00001111;
	mem[133] = 8'b00001111;
	mem[134] = 8'b00001111;
	mem[135] = 8'b00001111;
	mem[136] = 8'b00001111;
	mem[137] = 8'b00001111;
	mem[138] = 8'b00001111;
	mem[139] = 8'b00001111;
	mem[140] = 8'b00001101;
	mem[141] = 8'b00001010;
	mem[142] = 8'b00001010;
	mem[143] = 8'b00001010;
	mem[144] = 8'b00001010;
	mem[145] = 8'b00001010;
	mem[146] = 8'b00001010;
	mem[147] = 8'b00001010;
	mem[148] = 8'b00001010;
	mem[149] = 8'b00001010;
	mem[150] = 8'b00001010;
	mem[151] = 8'b00001010;
	mem[152] = 8'b00001010;
	mem[153] = 8'b00001010;
	mem[154] = 8'b00001010;
	mem[155] = 8'b00001011;
	mem[156] = 8'b00001111;
	mem[157] = 8'b00001111;
	mem[158] = 8'b00001111;
	mem[159] = 8'b00001111;
	mem[160] = 8'b00001111;
	mem[161] = 8'b00001111;
	mem[162] = 8'b00001111;
	mem[163] = 8'b00001111;
	mem[164] = 8'b00001111;
	mem[165] = 8'b00001111;
	mem[166] = 8'b00001111;
	mem[167] = 8'b00001111;
	mem[168] = 8'b00001111;
	mem[169] = 8'b00001111;
	mem[170] = 8'b00001111;
	mem[171] = 8'b00001111;
	mem[172] = 8'b00001111;
	mem[173] = 8'b00001111;
	mem[174] = 8'b00001111;
	mem[175] = 8'b00001111;
	mem[176] = 8'b00001111;
	mem[177] = 8'b00001111;
	mem[178] = 8'b00001111;
	mem[179] = 8'b00001111;
	mem[180] = 8'b00001111;
	mem[181] = 8'b00001111;
	mem[182] = 8'b00001111;
	mem[183] = 8'b00001111;
	mem[184] = 8'b00001111;
	mem[185] = 8'b00001111;
	mem[186] = 8'b00001111;
	mem[187] = 8'b00001111;
	mem[188] = 8'b00001111;
	mem[189] = 8'b00001111;
	mem[190] = 8'b00001111;
	mem[191] = 8'b00001111;
	mem[192] = 8'b00001111;
	mem[193] = 8'b00001111;
	mem[194] = 8'b00001111;
	mem[195] = 8'b00001111;
	mem[196] = 8'b00001111;
	mem[197] = 8'b00001111;
	mem[198] = 8'b00001111;
	mem[199] = 8'b00001111;
	mem[200] = 8'b00001111;
	mem[201] = 8'b00001111;
	mem[202] = 8'b00001111;
	mem[203] = 8'b00001100;
	mem[204] = 8'b00001010;
	mem[205] = 8'b00001010;
	mem[206] = 8'b00001010;
	mem[207] = 8'b00001010;
	mem[208] = 8'b00001010;
	mem[209] = 8'b00001010;
	mem[210] = 8'b00001011;
	mem[211] = 8'b00001011;
	mem[212] = 8'b00001011;
	mem[213] = 8'b00001011;
	mem[214] = 8'b00001010;
	mem[215] = 8'b00001010;
	mem[216] = 8'b00001010;
	mem[217] = 8'b00001010;
	mem[218] = 8'b00001010;
	mem[219] = 8'b00001010;
	mem[220] = 8'b00001111;
	mem[221] = 8'b00001111;
	mem[222] = 8'b00001111;
	mem[223] = 8'b00001111;
	mem[224] = 8'b00001111;
	mem[225] = 8'b00001111;
	mem[226] = 8'b00001111;
	mem[227] = 8'b00001111;
	mem[228] = 8'b00001111;
	mem[229] = 8'b00001111;
	mem[230] = 8'b00001111;
	mem[231] = 8'b00001111;
	mem[232] = 8'b00001111;
	mem[233] = 8'b00001111;
	mem[234] = 8'b00001111;
	mem[235] = 8'b00001111;
	mem[236] = 8'b00001111;
	mem[237] = 8'b00001111;
	mem[238] = 8'b00001111;
	mem[239] = 8'b00001111;
	mem[240] = 8'b00001111;
	mem[241] = 8'b00001111;
	mem[242] = 8'b00001111;
	mem[243] = 8'b00001111;
	mem[244] = 8'b00001111;
	mem[245] = 8'b00001111;
	mem[246] = 8'b00001111;
	mem[247] = 8'b00001111;
	mem[248] = 8'b00001111;
	mem[249] = 8'b00001111;
	mem[250] = 8'b00001111;
	mem[251] = 8'b00001111;
	mem[252] = 8'b00001111;
	mem[253] = 8'b00001111;
	mem[254] = 8'b00001111;
	mem[255] = 8'b00001111;
	mem[256] = 8'b00001111;
	mem[257] = 8'b00001111;
	mem[258] = 8'b00001111;
	mem[259] = 8'b00001111;
	mem[260] = 8'b00001101;
	mem[261] = 8'b00001011;
	mem[262] = 8'b00001010;
	mem[263] = 8'b00001011;
	mem[264] = 8'b00001011;
	mem[265] = 8'b00001011;
	mem[266] = 8'b00001011;
	mem[267] = 8'b00001010;
	mem[268] = 8'b00001010;
	mem[269] = 8'b00001010;
	mem[270] = 8'b00001010;
	mem[271] = 8'b00001010;
	mem[272] = 8'b00001011;
	mem[273] = 8'b00001100;
	mem[274] = 8'b00001100;
	mem[275] = 8'b00001100;
	mem[276] = 8'b00001100;
	mem[277] = 8'b00001100;
	mem[278] = 8'b00001100;
	mem[279] = 8'b00001100;
	mem[280] = 8'b00001011;
	mem[281] = 8'b00001010;
	mem[282] = 8'b00001010;
	mem[283] = 8'b00001010;
	mem[284] = 8'b00001011;
	mem[285] = 8'b00001010;
	mem[286] = 8'b00001010;
	mem[287] = 8'b00001010;
	mem[288] = 8'b00001010;
	mem[289] = 8'b00001010;
	mem[290] = 8'b00001011;
	mem[291] = 8'b00001111;
	mem[292] = 8'b00001100;
	mem[293] = 8'b00001010;
	mem[294] = 8'b00001010;
	mem[295] = 8'b00001010;
	mem[296] = 8'b00001010;
	mem[297] = 8'b00001011;
	mem[298] = 8'b00001110;
	mem[299] = 8'b00001111;
	mem[300] = 8'b00001111;
	mem[301] = 8'b00001100;
	mem[302] = 8'b00001010;
	mem[303] = 8'b00001010;
	mem[304] = 8'b00001010;
	mem[305] = 8'b00001011;
	mem[306] = 8'b00001110;
	mem[307] = 8'b00001110;
	mem[308] = 8'b00001011;
	mem[309] = 8'b00001010;
	mem[310] = 8'b00001010;
	mem[311] = 8'b00001010;
	mem[312] = 8'b00001010;
	mem[313] = 8'b00001010;
	mem[314] = 8'b00001010;
	mem[315] = 8'b00001011;
	mem[316] = 8'b00001011;
	mem[317] = 8'b00001100;
	mem[318] = 8'b00001111;
	mem[319] = 8'b00001111;
	mem[320] = 8'b00001111;
	mem[321] = 8'b00001111;
	mem[322] = 8'b00001111;
	mem[323] = 8'b00001011;
	mem[324] = 8'b00001010;
	mem[325] = 8'b00001010;
	mem[326] = 8'b00001010;
	mem[327] = 8'b00001010;
	mem[328] = 8'b00001010;
	mem[329] = 8'b00001010;
	mem[330] = 8'b00001010;
	mem[331] = 8'b00001010;
	mem[332] = 8'b00001010;
	mem[333] = 8'b00001010;
	mem[334] = 8'b00001011;
	mem[335] = 8'b00001100;
	mem[336] = 8'b00001100;
	mem[337] = 8'b00001100;
	mem[338] = 8'b00001100;
	mem[339] = 8'b00001100;
	mem[340] = 8'b00001100;
	mem[341] = 8'b00001100;
	mem[342] = 8'b00001100;
	mem[343] = 8'b00001100;
	mem[344] = 8'b00001010;
	mem[345] = 8'b00001010;
	mem[346] = 8'b00001010;
	mem[347] = 8'b00001010;
	mem[348] = 8'b00001010;
	mem[349] = 8'b00001010;
	mem[350] = 8'b00001010;
	mem[351] = 8'b00001010;
	mem[352] = 8'b00001010;
	mem[353] = 8'b00001010;
	mem[354] = 8'b00001010;
	mem[355] = 8'b00001010;
	mem[356] = 8'b00001010;
	mem[357] = 8'b00001010;
	mem[358] = 8'b00001010;
	mem[359] = 8'b00001010;
	mem[360] = 8'b00001010;
	mem[361] = 8'b00001010;
	mem[362] = 8'b00001010;
	mem[363] = 8'b00001101;
	mem[364] = 8'b00001011;
	mem[365] = 8'b00001010;
	mem[366] = 8'b00001010;
	mem[367] = 8'b00001010;
	mem[368] = 8'b00001010;
	mem[369] = 8'b00001010;
	mem[370] = 8'b00001010;
	mem[371] = 8'b00001010;
	mem[372] = 8'b00001010;
	mem[373] = 8'b00001010;
	mem[374] = 8'b00001010;
	mem[375] = 8'b00001010;
	mem[376] = 8'b00001010;
	mem[377] = 8'b00001010;
	mem[378] = 8'b00001010;
	mem[379] = 8'b00001010;
	mem[380] = 8'b00001010;
	mem[381] = 8'b00001010;
	mem[382] = 8'b00001010;
	mem[383] = 8'b00001111;
	mem[384] = 8'b00001111;
	mem[385] = 8'b00001111;
	mem[386] = 8'b00001110;
	mem[387] = 8'b00001010;
	mem[388] = 8'b00001010;
	mem[389] = 8'b00001010;
	mem[390] = 8'b00001010;
	mem[391] = 8'b00001010;
	mem[392] = 8'b00001010;
	mem[393] = 8'b00001010;
	mem[394] = 8'b00001010;
	mem[395] = 8'b00001010;
	mem[396] = 8'b00001010;
	mem[397] = 8'b00001011;
	mem[398] = 8'b00001100;
	mem[399] = 8'b00001100;
	mem[400] = 8'b00001100;
	mem[401] = 8'b00001011;
	mem[402] = 8'b00001011;
	mem[403] = 8'b00001010;
	mem[404] = 8'b00001011;
	mem[405] = 8'b00001011;
	mem[406] = 8'b00001100;
	mem[407] = 8'b00001011;
	mem[408] = 8'b00001010;
	mem[409] = 8'b00001010;
	mem[410] = 8'b00001010;
	mem[411] = 8'b00001010;
	mem[412] = 8'b00001010;
	mem[413] = 8'b00001010;
	mem[414] = 8'b00001010;
	mem[415] = 8'b00001010;
	mem[416] = 8'b00001010;
	mem[417] = 8'b00001010;
	mem[418] = 8'b00001010;
	mem[419] = 8'b00001010;
	mem[420] = 8'b00001010;
	mem[421] = 8'b00001010;
	mem[422] = 8'b00001010;
	mem[423] = 8'b00001010;
	mem[424] = 8'b00001010;
	mem[425] = 8'b00001010;
	mem[426] = 8'b00001010;
	mem[427] = 8'b00001010;
	mem[428] = 8'b00001010;
	mem[429] = 8'b00001010;
	mem[430] = 8'b00001010;
	mem[431] = 8'b00001010;
	mem[432] = 8'b00001010;
	mem[433] = 8'b00001010;
	mem[434] = 8'b00001010;
	mem[435] = 8'b00001010;
	mem[436] = 8'b00001010;
	mem[437] = 8'b00001010;
	mem[438] = 8'b00001010;
	mem[439] = 8'b00001010;
	mem[440] = 8'b00001010;
	mem[441] = 8'b00001010;
	mem[442] = 8'b00001010;
	mem[443] = 8'b00001010;
	mem[444] = 8'b00001010;
	mem[445] = 8'b00001010;
	mem[446] = 8'b00001010;
	mem[447] = 8'b00001011;
	mem[448] = 8'b00001111;
	mem[449] = 8'b00001111;
	mem[450] = 8'b00001011;
	mem[451] = 8'b00001010;
	mem[452] = 8'b00001010;
	mem[453] = 8'b00001010;
	mem[454] = 8'b00001010;
	mem[455] = 8'b00001010;
	mem[456] = 8'b00001010;
	mem[457] = 8'b00001010;
	mem[458] = 8'b00001010;
	mem[459] = 8'b00001010;
	mem[460] = 8'b00001100;
	mem[461] = 8'b00001100;
	mem[462] = 8'b00001100;
	mem[463] = 8'b00001100;
	mem[464] = 8'b00001010;
	mem[465] = 8'b00001010;
	mem[466] = 8'b00001010;
	mem[467] = 8'b00001010;
	mem[468] = 8'b00001010;
	mem[469] = 8'b00001010;
	mem[470] = 8'b00001010;
	mem[471] = 8'b00001010;
	mem[472] = 8'b00001010;
	mem[473] = 8'b00001010;
	mem[474] = 8'b00001010;
	mem[475] = 8'b00001010;
	mem[476] = 8'b00001010;
	mem[477] = 8'b00001010;
	mem[478] = 8'b00001010;
	mem[479] = 8'b00001010;
	mem[480] = 8'b00001010;
	mem[481] = 8'b00001010;
	mem[482] = 8'b00001010;
	mem[483] = 8'b00001010;
	mem[484] = 8'b00001010;
	mem[485] = 8'b00001010;
	mem[486] = 8'b00001010;
	mem[487] = 8'b00001010;
	mem[488] = 8'b00001010;
	mem[489] = 8'b00001010;
	mem[490] = 8'b00001010;
	mem[491] = 8'b00001010;
	mem[492] = 8'b00001010;
	mem[493] = 8'b00001010;
	mem[494] = 8'b00001010;
	mem[495] = 8'b00001010;
	mem[496] = 8'b00001010;
	mem[497] = 8'b00001010;
	mem[498] = 8'b00001010;
	mem[499] = 8'b00001010;
	mem[500] = 8'b00001010;
	mem[501] = 8'b00001010;
	mem[502] = 8'b00001010;
	mem[503] = 8'b00001010;
	mem[504] = 8'b00001010;
	mem[505] = 8'b00001010;
	mem[506] = 8'b00001010;
	mem[507] = 8'b00001010;
	mem[508] = 8'b00001010;
	mem[509] = 8'b00001010;
	mem[510] = 8'b00001010;
	mem[511] = 8'b00001010;
	mem[512] = 8'b00001111;
	mem[513] = 8'b00001111;
	mem[514] = 8'b00001011;
	mem[515] = 8'b00001010;
	mem[516] = 8'b00001010;
	mem[517] = 8'b00001010;
	mem[518] = 8'b00001100;
	mem[519] = 8'b00001100;
	mem[520] = 8'b00001100;
	mem[521] = 8'b00001100;
	mem[522] = 8'b00001100;
	mem[523] = 8'b00001100;
	mem[524] = 8'b00001100;
	mem[525] = 8'b00001100;
	mem[526] = 8'b00001100;
	mem[527] = 8'b00001010;
	mem[528] = 8'b00001010;
	mem[529] = 8'b00001100;
	mem[530] = 8'b00001011;
	mem[531] = 8'b00001010;
	mem[532] = 8'b00001010;
	mem[533] = 8'b00001010;
	mem[534] = 8'b00001010;
	mem[535] = 8'b00001010;
	mem[536] = 8'b00001010;
	mem[537] = 8'b00001010;
	mem[538] = 8'b00001010;
	mem[539] = 8'b00001010;
	mem[540] = 8'b00001010;
	mem[541] = 8'b00001011;
	mem[542] = 8'b00001100;
	mem[543] = 8'b00001100;
	mem[544] = 8'b00001100;
	mem[545] = 8'b00001010;
	mem[546] = 8'b00001010;
	mem[547] = 8'b00001010;
	mem[548] = 8'b00001010;
	mem[549] = 8'b00001010;
	mem[550] = 8'b00001100;
	mem[551] = 8'b00001100;
	mem[552] = 8'b00001011;
	mem[553] = 8'b00001010;
	mem[554] = 8'b00001010;
	mem[555] = 8'b00001010;
	mem[556] = 8'b00001010;
	mem[557] = 8'b00001010;
	mem[558] = 8'b00001011;
	mem[559] = 8'b00001100;
	mem[560] = 8'b00001100;
	mem[561] = 8'b00001011;
	mem[562] = 8'b00001010;
	mem[563] = 8'b00001010;
	mem[564] = 8'b00001010;
	mem[565] = 8'b00001100;
	mem[566] = 8'b00001100;
	mem[567] = 8'b00001100;
	mem[568] = 8'b00001100;
	mem[569] = 8'b00001100;
	mem[570] = 8'b00001100;
	mem[571] = 8'b00001100;
	mem[572] = 8'b00001010;
	mem[573] = 8'b00001010;
	mem[574] = 8'b00001010;
	mem[575] = 8'b00001010;
	mem[576] = 8'b00001111;
	mem[577] = 8'b00001111;
	mem[578] = 8'b00001100;
	mem[579] = 8'b00001010;
	mem[580] = 8'b00001010;
	mem[581] = 8'b00001010;
	mem[582] = 8'b00001100;
	mem[583] = 8'b00001100;
	mem[584] = 8'b00001100;
	mem[585] = 8'b00001100;
	mem[586] = 8'b00001100;
	mem[587] = 8'b00001100;
	mem[588] = 8'b00001100;
	mem[589] = 8'b00001011;
	mem[590] = 8'b00001010;
	mem[591] = 8'b00001010;
	mem[592] = 8'b00001011;
	mem[593] = 8'b00001100;
	mem[594] = 8'b00001100;
	mem[595] = 8'b00001010;
	mem[596] = 8'b00001010;
	mem[597] = 8'b00001010;
	mem[598] = 8'b00001010;
	mem[599] = 8'b00001010;
	mem[600] = 8'b00001010;
	mem[601] = 8'b00001010;
	mem[602] = 8'b00001010;
	mem[603] = 8'b00001010;
	mem[604] = 8'b00001010;
	mem[605] = 8'b00001100;
	mem[606] = 8'b00001100;
	mem[607] = 8'b00001100;
	mem[608] = 8'b00001100;
	mem[609] = 8'b00001010;
	mem[610] = 8'b00001010;
	mem[611] = 8'b00001010;
	mem[612] = 8'b00001010;
	mem[613] = 8'b00001011;
	mem[614] = 8'b00001100;
	mem[615] = 8'b00001100;
	mem[616] = 8'b00001100;
	mem[617] = 8'b00001011;
	mem[618] = 8'b00001010;
	mem[619] = 8'b00001010;
	mem[620] = 8'b00001010;
	mem[621] = 8'b00001100;
	mem[622] = 8'b00001100;
	mem[623] = 8'b00001100;
	mem[624] = 8'b00001100;
	mem[625] = 8'b00001011;
	mem[626] = 8'b00001010;
	mem[627] = 8'b00001010;
	mem[628] = 8'b00001010;
	mem[629] = 8'b00001100;
	mem[630] = 8'b00001100;
	mem[631] = 8'b00001100;
	mem[632] = 8'b00001100;
	mem[633] = 8'b00001100;
	mem[634] = 8'b00001100;
	mem[635] = 8'b00001100;
	mem[636] = 8'b00001010;
	mem[637] = 8'b00001010;
	mem[638] = 8'b00001010;
	mem[639] = 8'b00001010;
	mem[640] = 8'b00001111;
	mem[641] = 8'b00001111;
	mem[642] = 8'b00001011;
	mem[643] = 8'b00001001;
	mem[644] = 8'b00001001;
	mem[645] = 8'b00001001;
	mem[646] = 8'b00001100;
	mem[647] = 8'b00001100;
	mem[648] = 8'b00001100;
	mem[649] = 8'b00001011;
	mem[650] = 8'b00001011;
	mem[651] = 8'b00001010;
	mem[652] = 8'b00001010;
	mem[653] = 8'b00001001;
	mem[654] = 8'b00001001;
	mem[655] = 8'b00001001;
	mem[656] = 8'b00001011;
	mem[657] = 8'b00001100;
	mem[658] = 8'b00001100;
	mem[659] = 8'b00001001;
	mem[660] = 8'b00001001;
	mem[661] = 8'b00001001;
	mem[662] = 8'b00001010;
	mem[663] = 8'b00001011;
	mem[664] = 8'b00001001;
	mem[665] = 8'b00001001;
	mem[666] = 8'b00001001;
	mem[667] = 8'b00001010;
	mem[668] = 8'b00001100;
	mem[669] = 8'b00001100;
	mem[670] = 8'b00001100;
	mem[671] = 8'b00001100;
	mem[672] = 8'b00001100;
	mem[673] = 8'b00001001;
	mem[674] = 8'b00001001;
	mem[675] = 8'b00001001;
	mem[676] = 8'b00001001;
	mem[677] = 8'b00001100;
	mem[678] = 8'b00001100;
	mem[679] = 8'b00001100;
	mem[680] = 8'b00001100;
	mem[681] = 8'b00001100;
	mem[682] = 8'b00001010;
	mem[683] = 8'b00001010;
	mem[684] = 8'b00001100;
	mem[685] = 8'b00001100;
	mem[686] = 8'b00001100;
	mem[687] = 8'b00001100;
	mem[688] = 8'b00001100;
	mem[689] = 8'b00001010;
	mem[690] = 8'b00001001;
	mem[691] = 8'b00001001;
	mem[692] = 8'b00001011;
	mem[693] = 8'b00001100;
	mem[694] = 8'b00001100;
	mem[695] = 8'b00001011;
	mem[696] = 8'b00001011;
	mem[697] = 8'b00001011;
	mem[698] = 8'b00001011;
	mem[699] = 8'b00001011;
	mem[700] = 8'b00001010;
	mem[701] = 8'b00001001;
	mem[702] = 8'b00001001;
	mem[703] = 8'b00001010;
	mem[704] = 8'b00001111;
	mem[705] = 8'b00001111;
	mem[706] = 8'b00001010;
	mem[707] = 8'b00001001;
	mem[708] = 8'b00001001;
	mem[709] = 8'b00001010;
	mem[710] = 8'b00001100;
	mem[711] = 8'b00001100;
	mem[712] = 8'b00001010;
	mem[713] = 8'b00001001;
	mem[714] = 8'b00001001;
	mem[715] = 8'b00001001;
	mem[716] = 8'b00001001;
	mem[717] = 8'b00001001;
	mem[718] = 8'b00001001;
	mem[719] = 8'b00001001;
	mem[720] = 8'b00001100;
	mem[721] = 8'b00001100;
	mem[722] = 8'b00001011;
	mem[723] = 8'b00001001;
	mem[724] = 8'b00001001;
	mem[725] = 8'b00001001;
	mem[726] = 8'b00001011;
	mem[727] = 8'b00001010;
	mem[728] = 8'b00001001;
	mem[729] = 8'b00001001;
	mem[730] = 8'b00001001;
	mem[731] = 8'b00001011;
	mem[732] = 8'b00001100;
	mem[733] = 8'b00001100;
	mem[734] = 8'b00001100;
	mem[735] = 8'b00001100;
	mem[736] = 8'b00001100;
	mem[737] = 8'b00001010;
	mem[738] = 8'b00001001;
	mem[739] = 8'b00001001;
	mem[740] = 8'b00001010;
	mem[741] = 8'b00001100;
	mem[742] = 8'b00001100;
	mem[743] = 8'b00001100;
	mem[744] = 8'b00001100;
	mem[745] = 8'b00001100;
	mem[746] = 8'b00001100;
	mem[747] = 8'b00001100;
	mem[748] = 8'b00001100;
	mem[749] = 8'b00001100;
	mem[750] = 8'b00001100;
	mem[751] = 8'b00001100;
	mem[752] = 8'b00001100;
	mem[753] = 8'b00001001;
	mem[754] = 8'b00001001;
	mem[755] = 8'b00001001;
	mem[756] = 8'b00001100;
	mem[757] = 8'b00001100;
	mem[758] = 8'b00001100;
	mem[759] = 8'b00001001;
	mem[760] = 8'b00001001;
	mem[761] = 8'b00001001;
	mem[762] = 8'b00001001;
	mem[763] = 8'b00001001;
	mem[764] = 8'b00001001;
	mem[765] = 8'b00001001;
	mem[766] = 8'b00001001;
	mem[767] = 8'b00001010;
	mem[768] = 8'b00001111;
	mem[769] = 8'b00001111;
	mem[770] = 8'b00001001;
	mem[771] = 8'b00001001;
	mem[772] = 8'b00001001;
	mem[773] = 8'b00001011;
	mem[774] = 8'b00001100;
	mem[775] = 8'b00001100;
	mem[776] = 8'b00001011;
	mem[777] = 8'b00001010;
	mem[778] = 8'b00001010;
	mem[779] = 8'b00001010;
	mem[780] = 8'b00001001;
	mem[781] = 8'b00001001;
	mem[782] = 8'b00001001;
	mem[783] = 8'b00001010;
	mem[784] = 8'b00001100;
	mem[785] = 8'b00001100;
	mem[786] = 8'b00001010;
	mem[787] = 8'b00001001;
	mem[788] = 8'b00001001;
	mem[789] = 8'b00001001;
	mem[790] = 8'b00001010;
	mem[791] = 8'b00001001;
	mem[792] = 8'b00001001;
	mem[793] = 8'b00001001;
	mem[794] = 8'b00001010;
	mem[795] = 8'b00001100;
	mem[796] = 8'b00001100;
	mem[797] = 8'b00001100;
	mem[798] = 8'b00001010;
	mem[799] = 8'b00001100;
	mem[800] = 8'b00001100;
	mem[801] = 8'b00001010;
	mem[802] = 8'b00001001;
	mem[803] = 8'b00001001;
	mem[804] = 8'b00001010;
	mem[805] = 8'b00001100;
	mem[806] = 8'b00001100;
	mem[807] = 8'b00001010;
	mem[808] = 8'b00001011;
	mem[809] = 8'b00001100;
	mem[810] = 8'b00001100;
	mem[811] = 8'b00001100;
	mem[812] = 8'b00001100;
	mem[813] = 8'b00001011;
	mem[814] = 8'b00001100;
	mem[815] = 8'b00001100;
	mem[816] = 8'b00001011;
	mem[817] = 8'b00001001;
	mem[818] = 8'b00001001;
	mem[819] = 8'b00001001;
	mem[820] = 8'b00001100;
	mem[821] = 8'b00001100;
	mem[822] = 8'b00001100;
	mem[823] = 8'b00001011;
	mem[824] = 8'b00001011;
	mem[825] = 8'b00001011;
	mem[826] = 8'b00001010;
	mem[827] = 8'b00001001;
	mem[828] = 8'b00001001;
	mem[829] = 8'b00001001;
	mem[830] = 8'b00001001;
	mem[831] = 8'b00001101;
	mem[832] = 8'b00001111;
	mem[833] = 8'b00001100;
	mem[834] = 8'b00001001;
	mem[835] = 8'b00001001;
	mem[836] = 8'b00001001;
	mem[837] = 8'b00001100;
	mem[838] = 8'b00001100;
	mem[839] = 8'b00001100;
	mem[840] = 8'b00001100;
	mem[841] = 8'b00001100;
	mem[842] = 8'b00001100;
	mem[843] = 8'b00001100;
	mem[844] = 8'b00001001;
	mem[845] = 8'b00001001;
	mem[846] = 8'b00001001;
	mem[847] = 8'b00001011;
	mem[848] = 8'b00001100;
	mem[849] = 8'b00001100;
	mem[850] = 8'b00001001;
	mem[851] = 8'b00001001;
	mem[852] = 8'b00001001;
	mem[853] = 8'b00001001;
	mem[854] = 8'b00001001;
	mem[855] = 8'b00001001;
	mem[856] = 8'b00001001;
	mem[857] = 8'b00001001;
	mem[858] = 8'b00001100;
	mem[859] = 8'b00001100;
	mem[860] = 8'b00001100;
	mem[861] = 8'b00001010;
	mem[862] = 8'b00001001;
	mem[863] = 8'b00001100;
	mem[864] = 8'b00001100;
	mem[865] = 8'b00001010;
	mem[866] = 8'b00001001;
	mem[867] = 8'b00001001;
	mem[868] = 8'b00001011;
	mem[869] = 8'b00001100;
	mem[870] = 8'b00001100;
	mem[871] = 8'b00001001;
	mem[872] = 8'b00001001;
	mem[873] = 8'b00001100;
	mem[874] = 8'b00001100;
	mem[875] = 8'b00001100;
	mem[876] = 8'b00001001;
	mem[877] = 8'b00001010;
	mem[878] = 8'b00001100;
	mem[879] = 8'b00001100;
	mem[880] = 8'b00001010;
	mem[881] = 8'b00001001;
	mem[882] = 8'b00001001;
	mem[883] = 8'b00001010;
	mem[884] = 8'b00001100;
	mem[885] = 8'b00001100;
	mem[886] = 8'b00001100;
	mem[887] = 8'b00001100;
	mem[888] = 8'b00001100;
	mem[889] = 8'b00001100;
	mem[890] = 8'b00001010;
	mem[891] = 8'b00001001;
	mem[892] = 8'b00001001;
	mem[893] = 8'b00001001;
	mem[894] = 8'b00001100;
	mem[895] = 8'b00001111;
	mem[896] = 8'b00001111;
	mem[897] = 8'b00001010;
	mem[898] = 8'b00001001;
	mem[899] = 8'b00001001;
	mem[900] = 8'b00001001;
	mem[901] = 8'b00001100;
	mem[902] = 8'b00001100;
	mem[903] = 8'b00001100;
	mem[904] = 8'b00001100;
	mem[905] = 8'b00001100;
	mem[906] = 8'b00001100;
	mem[907] = 8'b00001100;
	mem[908] = 8'b00001001;
	mem[909] = 8'b00001001;
	mem[910] = 8'b00001001;
	mem[911] = 8'b00001100;
	mem[912] = 8'b00001100;
	mem[913] = 8'b00001100;
	mem[914] = 8'b00001001;
	mem[915] = 8'b00001001;
	mem[916] = 8'b00001001;
	mem[917] = 8'b00001001;
	mem[918] = 8'b00001001;
	mem[919] = 8'b00001001;
	mem[920] = 8'b00001001;
	mem[921] = 8'b00001011;
	mem[922] = 8'b00001100;
	mem[923] = 8'b00001100;
	mem[924] = 8'b00001011;
	mem[925] = 8'b00001001;
	mem[926] = 8'b00001001;
	mem[927] = 8'b00001100;
	mem[928] = 8'b00001100;
	mem[929] = 8'b00001011;
	mem[930] = 8'b00001001;
	mem[931] = 8'b00001001;
	mem[932] = 8'b00001100;
	mem[933] = 8'b00001100;
	mem[934] = 8'b00001011;
	mem[935] = 8'b00001001;
	mem[936] = 8'b00001001;
	mem[937] = 8'b00001010;
	mem[938] = 8'b00001011;
	mem[939] = 8'b00001001;
	mem[940] = 8'b00001001;
	mem[941] = 8'b00001011;
	mem[942] = 8'b00001100;
	mem[943] = 8'b00001100;
	mem[944] = 8'b00001001;
	mem[945] = 8'b00001001;
	mem[946] = 8'b00001001;
	mem[947] = 8'b00001011;
	mem[948] = 8'b00001100;
	mem[949] = 8'b00001100;
	mem[950] = 8'b00001100;
	mem[951] = 8'b00001100;
	mem[952] = 8'b00001100;
	mem[953] = 8'b00001100;
	mem[954] = 8'b00001010;
	mem[955] = 8'b00001001;
	mem[956] = 8'b00001001;
	mem[957] = 8'b00001001;
	mem[958] = 8'b00001111;
	mem[959] = 8'b00001111;
	mem[960] = 8'b00001111;
	mem[961] = 8'b00001001;
	mem[962] = 8'b00001001;
	mem[963] = 8'b00001001;
	mem[964] = 8'b00001010;
	mem[965] = 8'b00001100;
	mem[966] = 8'b00001100;
	mem[967] = 8'b00001010;
	mem[968] = 8'b00001001;
	mem[969] = 8'b00001001;
	mem[970] = 8'b00001001;
	mem[971] = 8'b00001001;
	mem[972] = 8'b00001001;
	mem[973] = 8'b00001001;
	mem[974] = 8'b00001001;
	mem[975] = 8'b00001100;
	mem[976] = 8'b00001100;
	mem[977] = 8'b00001011;
	mem[978] = 8'b00001001;
	mem[979] = 8'b00001001;
	mem[980] = 8'b00001001;
	mem[981] = 8'b00001001;
	mem[982] = 8'b00001001;
	mem[983] = 8'b00001001;
	mem[984] = 8'b00001010;
	mem[985] = 8'b00001100;
	mem[986] = 8'b00001100;
	mem[987] = 8'b00001100;
	mem[988] = 8'b00001100;
	mem[989] = 8'b00001100;
	mem[990] = 8'b00001100;
	mem[991] = 8'b00001100;
	mem[992] = 8'b00001100;
	mem[993] = 8'b00001011;
	mem[994] = 8'b00001001;
	mem[995] = 8'b00001010;
	mem[996] = 8'b00001100;
	mem[997] = 8'b00001100;
	mem[998] = 8'b00001010;
	mem[999] = 8'b00001001;
	mem[1000] = 8'b00001001;
	mem[1001] = 8'b00001001;
	mem[1002] = 8'b00001001;
	mem[1003] = 8'b00001001;
	mem[1004] = 8'b00001001;
	mem[1005] = 8'b00001100;
	mem[1006] = 8'b00001100;
	mem[1007] = 8'b00001011;
	mem[1008] = 8'b00001001;
	mem[1009] = 8'b00001001;
	mem[1010] = 8'b00001001;
	mem[1011] = 8'b00001100;
	mem[1012] = 8'b00001100;
	mem[1013] = 8'b00001011;
	mem[1014] = 8'b00001001;
	mem[1015] = 8'b00001001;
	mem[1016] = 8'b00001001;
	mem[1017] = 8'b00001001;
	mem[1018] = 8'b00001001;
	mem[1019] = 8'b00001001;
	mem[1020] = 8'b00001001;
	mem[1021] = 8'b00001001;
	mem[1022] = 8'b00001111;
	mem[1023] = 8'b00001111;
	mem[1024] = 8'b00001101;
	mem[1025] = 8'b00001001;
	mem[1026] = 8'b00001001;
	mem[1027] = 8'b00001001;
	mem[1028] = 8'b00001011;
	mem[1029] = 8'b00001100;
	mem[1030] = 8'b00001100;
	mem[1031] = 8'b00001001;
	mem[1032] = 8'b00001001;
	mem[1033] = 8'b00001001;
	mem[1034] = 8'b00001001;
	mem[1035] = 8'b00001001;
	mem[1036] = 8'b00001001;
	mem[1037] = 8'b00001001;
	mem[1038] = 8'b00001010;
	mem[1039] = 8'b00001100;
	mem[1040] = 8'b00001100;
	mem[1041] = 8'b00001001;
	mem[1042] = 8'b00001001;
	mem[1043] = 8'b00001001;
	mem[1044] = 8'b00001001;
	mem[1045] = 8'b00001001;
	mem[1046] = 8'b00001001;
	mem[1047] = 8'b00001001;
	mem[1048] = 8'b00001100;
	mem[1049] = 8'b00001100;
	mem[1050] = 8'b00001100;
	mem[1051] = 8'b00001100;
	mem[1052] = 8'b00001100;
	mem[1053] = 8'b00001100;
	mem[1054] = 8'b00001100;
	mem[1055] = 8'b00001100;
	mem[1056] = 8'b00001100;
	mem[1057] = 8'b00001011;
	mem[1058] = 8'b00001001;
	mem[1059] = 8'b00001011;
	mem[1060] = 8'b00001100;
	mem[1061] = 8'b00001100;
	mem[1062] = 8'b00001001;
	mem[1063] = 8'b00001001;
	mem[1064] = 8'b00001001;
	mem[1065] = 8'b00001001;
	mem[1066] = 8'b00001001;
	mem[1067] = 8'b00001001;
	mem[1068] = 8'b00001010;
	mem[1069] = 8'b00001100;
	mem[1070] = 8'b00001100;
	mem[1071] = 8'b00001010;
	mem[1072] = 8'b00001001;
	mem[1073] = 8'b00001001;
	mem[1074] = 8'b00001001;
	mem[1075] = 8'b00001100;
	mem[1076] = 8'b00001100;
	mem[1077] = 8'b00001010;
	mem[1078] = 8'b00001001;
	mem[1079] = 8'b00001001;
	mem[1080] = 8'b00001001;
	mem[1081] = 8'b00001001;
	mem[1082] = 8'b00001001;
	mem[1083] = 8'b00001001;
	mem[1084] = 8'b00001001;
	mem[1085] = 8'b00001010;
	mem[1086] = 8'b00001111;
	mem[1087] = 8'b00001111;
	mem[1088] = 8'b00001010;
	mem[1089] = 8'b00001000;
	mem[1090] = 8'b00001000;
	mem[1091] = 8'b00001001;
	mem[1092] = 8'b00001100;
	mem[1093] = 8'b00001100;
	mem[1094] = 8'b00001011;
	mem[1095] = 8'b00001000;
	mem[1096] = 8'b00001000;
	mem[1097] = 8'b00001000;
	mem[1098] = 8'b00001000;
	mem[1099] = 8'b00001000;
	mem[1100] = 8'b00001000;
	mem[1101] = 8'b00001000;
	mem[1102] = 8'b00001011;
	mem[1103] = 8'b00001100;
	mem[1104] = 8'b00001100;
	mem[1105] = 8'b00001011;
	mem[1106] = 8'b00001011;
	mem[1107] = 8'b00001011;
	mem[1108] = 8'b00001011;
	mem[1109] = 8'b00001011;
	mem[1110] = 8'b00001001;
	mem[1111] = 8'b00001011;
	mem[1112] = 8'b00001100;
	mem[1113] = 8'b00001100;
	mem[1114] = 8'b00001011;
	mem[1115] = 8'b00001010;
	mem[1116] = 8'b00001010;
	mem[1117] = 8'b00001010;
	mem[1118] = 8'b00001010;
	mem[1119] = 8'b00001100;
	mem[1120] = 8'b00001100;
	mem[1121] = 8'b00001100;
	mem[1122] = 8'b00001000;
	mem[1123] = 8'b00001100;
	mem[1124] = 8'b00001100;
	mem[1125] = 8'b00001100;
	mem[1126] = 8'b00001000;
	mem[1127] = 8'b00001000;
	mem[1128] = 8'b00001000;
	mem[1129] = 8'b00001000;
	mem[1130] = 8'b00001000;
	mem[1131] = 8'b00001000;
	mem[1132] = 8'b00001011;
	mem[1133] = 8'b00001100;
	mem[1134] = 8'b00001100;
	mem[1135] = 8'b00001001;
	mem[1136] = 8'b00001000;
	mem[1137] = 8'b00001000;
	mem[1138] = 8'b00001010;
	mem[1139] = 8'b00001100;
	mem[1140] = 8'b00001100;
	mem[1141] = 8'b00001100;
	mem[1142] = 8'b00001100;
	mem[1143] = 8'b00001100;
	mem[1144] = 8'b00001100;
	mem[1145] = 8'b00001011;
	mem[1146] = 8'b00001000;
	mem[1147] = 8'b00001000;
	mem[1148] = 8'b00001000;
	mem[1149] = 8'b00001010;
	mem[1150] = 8'b00001111;
	mem[1151] = 8'b00001111;
	mem[1152] = 8'b00001001;
	mem[1153] = 8'b00001000;
	mem[1154] = 8'b00001000;
	mem[1155] = 8'b00001001;
	mem[1156] = 8'b00001100;
	mem[1157] = 8'b00001100;
	mem[1158] = 8'b00001010;
	mem[1159] = 8'b00001000;
	mem[1160] = 8'b00001000;
	mem[1161] = 8'b00001000;
	mem[1162] = 8'b00001001;
	mem[1163] = 8'b00001000;
	mem[1164] = 8'b00001000;
	mem[1165] = 8'b00001000;
	mem[1166] = 8'b00001100;
	mem[1167] = 8'b00001100;
	mem[1168] = 8'b00001100;
	mem[1169] = 8'b00001100;
	mem[1170] = 8'b00001100;
	mem[1171] = 8'b00001100;
	mem[1172] = 8'b00001100;
	mem[1173] = 8'b00001100;
	mem[1174] = 8'b00001010;
	mem[1175] = 8'b00001100;
	mem[1176] = 8'b00001100;
	mem[1177] = 8'b00001011;
	mem[1178] = 8'b00001000;
	mem[1179] = 8'b00001000;
	mem[1180] = 8'b00001000;
	mem[1181] = 8'b00001000;
	mem[1182] = 8'b00001000;
	mem[1183] = 8'b00001010;
	mem[1184] = 8'b00001100;
	mem[1185] = 8'b00001100;
	mem[1186] = 8'b00001001;
	mem[1187] = 8'b00001100;
	mem[1188] = 8'b00001100;
	mem[1189] = 8'b00001010;
	mem[1190] = 8'b00001000;
	mem[1191] = 8'b00001000;
	mem[1192] = 8'b00001000;
	mem[1193] = 8'b00001000;
	mem[1194] = 8'b00001000;
	mem[1195] = 8'b00001000;
	mem[1196] = 8'b00001100;
	mem[1197] = 8'b00001100;
	mem[1198] = 8'b00001100;
	mem[1199] = 8'b00001000;
	mem[1200] = 8'b00001000;
	mem[1201] = 8'b00001000;
	mem[1202] = 8'b00001100;
	mem[1203] = 8'b00001100;
	mem[1204] = 8'b00001100;
	mem[1205] = 8'b00001100;
	mem[1206] = 8'b00001100;
	mem[1207] = 8'b00001100;
	mem[1208] = 8'b00001100;
	mem[1209] = 8'b00001100;
	mem[1210] = 8'b00001000;
	mem[1211] = 8'b00001000;
	mem[1212] = 8'b00001000;
	mem[1213] = 8'b00001010;
	mem[1214] = 8'b00001111;
	mem[1215] = 8'b00001111;
	mem[1216] = 8'b00001001;
	mem[1217] = 8'b00001000;
	mem[1218] = 8'b00001000;
	mem[1219] = 8'b00001001;
	mem[1220] = 8'b00001100;
	mem[1221] = 8'b00001100;
	mem[1222] = 8'b00001001;
	mem[1223] = 8'b00001000;
	mem[1224] = 8'b00001000;
	mem[1225] = 8'b00001000;
	mem[1226] = 8'b00001010;
	mem[1227] = 8'b00001000;
	mem[1228] = 8'b00001000;
	mem[1229] = 8'b00001001;
	mem[1230] = 8'b00001011;
	mem[1231] = 8'b00001100;
	mem[1232] = 8'b00001100;
	mem[1233] = 8'b00001100;
	mem[1234] = 8'b00001100;
	mem[1235] = 8'b00001100;
	mem[1236] = 8'b00001100;
	mem[1237] = 8'b00001100;
	mem[1238] = 8'b00001001;
	mem[1239] = 8'b00001011;
	mem[1240] = 8'b00001100;
	mem[1241] = 8'b00001001;
	mem[1242] = 8'b00001000;
	mem[1243] = 8'b00001000;
	mem[1244] = 8'b00001000;
	mem[1245] = 8'b00001000;
	mem[1246] = 8'b00001000;
	mem[1247] = 8'b00001010;
	mem[1248] = 8'b00001011;
	mem[1249] = 8'b00001011;
	mem[1250] = 8'b00001001;
	mem[1251] = 8'b00001011;
	mem[1252] = 8'b00001100;
	mem[1253] = 8'b00001001;
	mem[1254] = 8'b00001000;
	mem[1255] = 8'b00001000;
	mem[1256] = 8'b00001000;
	mem[1257] = 8'b00001000;
	mem[1258] = 8'b00001000;
	mem[1259] = 8'b00001000;
	mem[1260] = 8'b00001011;
	mem[1261] = 8'b00001011;
	mem[1262] = 8'b00001010;
	mem[1263] = 8'b00001000;
	mem[1264] = 8'b00001000;
	mem[1265] = 8'b00001000;
	mem[1266] = 8'b00001010;
	mem[1267] = 8'b00001100;
	mem[1268] = 8'b00001011;
	mem[1269] = 8'b00001011;
	mem[1270] = 8'b00001011;
	mem[1271] = 8'b00001011;
	mem[1272] = 8'b00001011;
	mem[1273] = 8'b00001011;
	mem[1274] = 8'b00001000;
	mem[1275] = 8'b00001000;
	mem[1276] = 8'b00001000;
	mem[1277] = 8'b00001010;
	mem[1278] = 8'b00001111;
	mem[1279] = 8'b00001111;
	mem[1280] = 8'b00001010;
	mem[1281] = 8'b00001000;
	mem[1282] = 8'b00001000;
	mem[1283] = 8'b00001000;
	mem[1284] = 8'b00001000;
	mem[1285] = 8'b00001001;
	mem[1286] = 8'b00001000;
	mem[1287] = 8'b00001000;
	mem[1288] = 8'b00001000;
	mem[1289] = 8'b00001001;
	mem[1290] = 8'b00001011;
	mem[1291] = 8'b00001000;
	mem[1292] = 8'b00001000;
	mem[1293] = 8'b00001000;
	mem[1294] = 8'b00001000;
	mem[1295] = 8'b00001000;
	mem[1296] = 8'b00001000;
	mem[1297] = 8'b00001000;
	mem[1298] = 8'b00001000;
	mem[1299] = 8'b00001000;
	mem[1300] = 8'b00001000;
	mem[1301] = 8'b00001000;
	mem[1302] = 8'b00001000;
	mem[1303] = 8'b00001000;
	mem[1304] = 8'b00001001;
	mem[1305] = 8'b00001000;
	mem[1306] = 8'b00001000;
	mem[1307] = 8'b00001000;
	mem[1308] = 8'b00001000;
	mem[1309] = 8'b00001000;
	mem[1310] = 8'b00001000;
	mem[1311] = 8'b00001000;
	mem[1312] = 8'b00001000;
	mem[1313] = 8'b00001000;
	mem[1314] = 8'b00001000;
	mem[1315] = 8'b00001000;
	mem[1316] = 8'b00001000;
	mem[1317] = 8'b00001000;
	mem[1318] = 8'b00001000;
	mem[1319] = 8'b00001000;
	mem[1320] = 8'b00001000;
	mem[1321] = 8'b00001000;
	mem[1322] = 8'b00001000;
	mem[1323] = 8'b00001000;
	mem[1324] = 8'b00001000;
	mem[1325] = 8'b00001000;
	mem[1326] = 8'b00001000;
	mem[1327] = 8'b00001000;
	mem[1328] = 8'b00001000;
	mem[1329] = 8'b00001000;
	mem[1330] = 8'b00001000;
	mem[1331] = 8'b00001000;
	mem[1332] = 8'b00001000;
	mem[1333] = 8'b00001000;
	mem[1334] = 8'b00001000;
	mem[1335] = 8'b00001000;
	mem[1336] = 8'b00001000;
	mem[1337] = 8'b00001000;
	mem[1338] = 8'b00001000;
	mem[1339] = 8'b00001000;
	mem[1340] = 8'b00001000;
	mem[1341] = 8'b00001011;
	mem[1342] = 8'b00001111;
	mem[1343] = 8'b00001111;
	mem[1344] = 8'b00001100;
	mem[1345] = 8'b00001000;
	mem[1346] = 8'b00001000;
	mem[1347] = 8'b00001000;
	mem[1348] = 8'b00001000;
	mem[1349] = 8'b00001000;
	mem[1350] = 8'b00001000;
	mem[1351] = 8'b00001000;
	mem[1352] = 8'b00001000;
	mem[1353] = 8'b00001011;
	mem[1354] = 8'b00001111;
	mem[1355] = 8'b00001001;
	mem[1356] = 8'b00001000;
	mem[1357] = 8'b00001000;
	mem[1358] = 8'b00001000;
	mem[1359] = 8'b00001000;
	mem[1360] = 8'b00001000;
	mem[1361] = 8'b00001000;
	mem[1362] = 8'b00001000;
	mem[1363] = 8'b00001000;
	mem[1364] = 8'b00001000;
	mem[1365] = 8'b00001000;
	mem[1366] = 8'b00001000;
	mem[1367] = 8'b00001000;
	mem[1368] = 8'b00001000;
	mem[1369] = 8'b00001000;
	mem[1370] = 8'b00001000;
	mem[1371] = 8'b00001000;
	mem[1372] = 8'b00001010;
	mem[1373] = 8'b00001000;
	mem[1374] = 8'b00001000;
	mem[1375] = 8'b00001000;
	mem[1376] = 8'b00001000;
	mem[1377] = 8'b00001000;
	mem[1378] = 8'b00001000;
	mem[1379] = 8'b00001000;
	mem[1380] = 8'b00001000;
	mem[1381] = 8'b00001000;
	mem[1382] = 8'b00001000;
	mem[1383] = 8'b00001000;
	mem[1384] = 8'b00001010;
	mem[1385] = 8'b00001001;
	mem[1386] = 8'b00001000;
	mem[1387] = 8'b00001000;
	mem[1388] = 8'b00001000;
	mem[1389] = 8'b00001000;
	mem[1390] = 8'b00001000;
	mem[1391] = 8'b00001000;
	mem[1392] = 8'b00001000;
	mem[1393] = 8'b00001000;
	mem[1394] = 8'b00001000;
	mem[1395] = 8'b00001000;
	mem[1396] = 8'b00001000;
	mem[1397] = 8'b00001000;
	mem[1398] = 8'b00001000;
	mem[1399] = 8'b00001000;
	mem[1400] = 8'b00001000;
	mem[1401] = 8'b00001000;
	mem[1402] = 8'b00001000;
	mem[1403] = 8'b00001000;
	mem[1404] = 8'b00001000;
	mem[1405] = 8'b00001110;
	mem[1406] = 8'b00001111;
	mem[1407] = 8'b00001111;
	mem[1408] = 8'b00001111;
	mem[1409] = 8'b00001100;
	mem[1410] = 8'b00001001;
	mem[1411] = 8'b00001000;
	mem[1412] = 8'b00001000;
	mem[1413] = 8'b00001000;
	mem[1414] = 8'b00001000;
	mem[1415] = 8'b00001000;
	mem[1416] = 8'b00001001;
	mem[1417] = 8'b00001111;
	mem[1418] = 8'b00001111;
	mem[1419] = 8'b00001110;
	mem[1420] = 8'b00001010;
	mem[1421] = 8'b00001000;
	mem[1422] = 8'b00001000;
	mem[1423] = 8'b00001000;
	mem[1424] = 8'b00001000;
	mem[1425] = 8'b00001000;
	mem[1426] = 8'b00001000;
	mem[1427] = 8'b00001000;
	mem[1428] = 8'b00001000;
	mem[1429] = 8'b00001000;
	mem[1430] = 8'b00001000;
	mem[1431] = 8'b00001000;
	mem[1432] = 8'b00001000;
	mem[1433] = 8'b00001000;
	mem[1434] = 8'b00001000;
	mem[1435] = 8'b00001011;
	mem[1436] = 8'b00001111;
	mem[1437] = 8'b00001010;
	mem[1438] = 8'b00001000;
	mem[1439] = 8'b00001000;
	mem[1440] = 8'b00001000;
	mem[1441] = 8'b00001000;
	mem[1442] = 8'b00001000;
	mem[1443] = 8'b00001000;
	mem[1444] = 8'b00001000;
	mem[1445] = 8'b00001000;
	mem[1446] = 8'b00001000;
	mem[1447] = 8'b00001001;
	mem[1448] = 8'b00001111;
	mem[1449] = 8'b00001101;
	mem[1450] = 8'b00001001;
	mem[1451] = 8'b00001000;
	mem[1452] = 8'b00001000;
	mem[1453] = 8'b00001000;
	mem[1454] = 8'b00001000;
	mem[1455] = 8'b00001000;
	mem[1456] = 8'b00001001;
	mem[1457] = 8'b00001001;
	mem[1458] = 8'b00001000;
	mem[1459] = 8'b00001000;
	mem[1460] = 8'b00001000;
	mem[1461] = 8'b00001000;
	mem[1462] = 8'b00001000;
	mem[1463] = 8'b00001000;
	mem[1464] = 8'b00001000;
	mem[1465] = 8'b00001000;
	mem[1466] = 8'b00001000;
	mem[1467] = 8'b00001001;
	mem[1468] = 8'b00001100;
	mem[1469] = 8'b00001111;
	mem[1470] = 8'b00001111;
	mem[1471] = 8'b00001111;
	mem[1472] = 8'b00001111;
	mem[1473] = 8'b00001111;
	mem[1474] = 8'b00001111;
	mem[1475] = 8'b00001101;
	mem[1476] = 8'b00001010;
	mem[1477] = 8'b00001001;
	mem[1478] = 8'b00001001;
	mem[1479] = 8'b00001011;
	mem[1480] = 8'b00001111;
	mem[1481] = 8'b00001111;
	mem[1482] = 8'b00001111;
	mem[1483] = 8'b00001111;
	mem[1484] = 8'b00001111;
	mem[1485] = 8'b00001110;
	mem[1486] = 8'b00001011;
	mem[1487] = 8'b00001001;
	mem[1488] = 8'b00001001;
	mem[1489] = 8'b00001010;
	mem[1490] = 8'b00001010;
	mem[1491] = 8'b00001010;
	mem[1492] = 8'b00001010;
	mem[1493] = 8'b00001010;
	mem[1494] = 8'b00001010;
	mem[1495] = 8'b00001001;
	mem[1496] = 8'b00001001;
	mem[1497] = 8'b00001001;
	mem[1498] = 8'b00001100;
	mem[1499] = 8'b00001111;
	mem[1500] = 8'b00001111;
	mem[1501] = 8'b00001111;
	mem[1502] = 8'b00001110;
	mem[1503] = 8'b00001011;
	mem[1504] = 8'b00001011;
	mem[1505] = 8'b00001100;
	mem[1506] = 8'b00001011;
	mem[1507] = 8'b00001011;
	mem[1508] = 8'b00001010;
	mem[1509] = 8'b00001010;
	mem[1510] = 8'b00001100;
	mem[1511] = 8'b00001111;
	mem[1512] = 8'b00001111;
	mem[1513] = 8'b00001111;
	mem[1514] = 8'b00001111;
	mem[1515] = 8'b00001101;
	mem[1516] = 8'b00001011;
	mem[1517] = 8'b00001010;
	mem[1518] = 8'b00001010;
	mem[1519] = 8'b00001011;
	mem[1520] = 8'b00001111;
	mem[1521] = 8'b00001111;
	mem[1522] = 8'b00001101;
	mem[1523] = 8'b00001010;
	mem[1524] = 8'b00001010;
	mem[1525] = 8'b00001011;
	mem[1526] = 8'b00001110;
	mem[1527] = 8'b00001111;
	mem[1528] = 8'b00001101;
	mem[1529] = 8'b00001011;
	mem[1530] = 8'b00001100;
	mem[1531] = 8'b00001111;
	mem[1532] = 8'b00001111;
	mem[1533] = 8'b00001111;
	mem[1534] = 8'b00001111;
	mem[1535] = 8'b00001111;
	mem[1536] = 8'b00000000;
	mem[1537] = 8'b00000000;
	mem[1538] = 8'b00000000;
	mem[1539] = 8'b00000000;
	mem[1540] = 8'b00000000;
	mem[1541] = 8'b00000000;
	mem[1542] = 8'b00000000;
	mem[1543] = 8'b00000000;
	mem[1544] = 8'b00000000;
	mem[1545] = 8'b00000000;
	mem[1546] = 8'b00000000;
	mem[1547] = 8'b00000000;
	mem[1548] = 8'b00000000;
	mem[1549] = 8'b00000000;
	mem[1550] = 8'b00000000;
	mem[1551] = 8'b00000000;
	mem[1552] = 8'b00000000;
	mem[1553] = 8'b00000000;
	mem[1554] = 8'b00000000;
	mem[1555] = 8'b00000000;
	mem[1556] = 8'b00000000;
	mem[1557] = 8'b00000000;
	mem[1558] = 8'b00000000;
	mem[1559] = 8'b00000000;
	mem[1560] = 8'b00000000;
	mem[1561] = 8'b00000000;
	mem[1562] = 8'b00000000;
	mem[1563] = 8'b00000000;
	mem[1564] = 8'b00000000;
	mem[1565] = 8'b00000000;
	mem[1566] = 8'b00000000;
	mem[1567] = 8'b00000000;
	mem[1568] = 8'b00000000;
	mem[1569] = 8'b00000000;
	mem[1570] = 8'b00000000;
	mem[1571] = 8'b00000000;
	mem[1572] = 8'b00000000;
	mem[1573] = 8'b00000000;
	mem[1574] = 8'b00000000;
	mem[1575] = 8'b00000000;
	mem[1576] = 8'b00000000;
	mem[1577] = 8'b00000000;
	mem[1578] = 8'b00000000;
	mem[1579] = 8'b00000000;
	mem[1580] = 8'b00000000;
	mem[1581] = 8'b00000000;
	mem[1582] = 8'b00000000;
	mem[1583] = 8'b00000000;
	mem[1584] = 8'b00000000;
	mem[1585] = 8'b00000000;
	mem[1586] = 8'b00000000;
	mem[1587] = 8'b00000000;
	mem[1588] = 8'b00000000;
	mem[1589] = 8'b00000000;
	mem[1590] = 8'b00000000;
	mem[1591] = 8'b00000000;
	mem[1592] = 8'b00000000;
	mem[1593] = 8'b00000000;
	mem[1594] = 8'b00000000;
	mem[1595] = 8'b00000000;
	mem[1596] = 8'b00000000;
	mem[1597] = 8'b00000000;
	mem[1598] = 8'b00000000;
	mem[1599] = 8'b00000000;
	mem[1600] = 8'b00000000;
	mem[1601] = 8'b00000000;
	mem[1602] = 8'b00000000;
	mem[1603] = 8'b00000000;
	mem[1604] = 8'b00000000;
	mem[1605] = 8'b00000000;
	mem[1606] = 8'b00000000;
	mem[1607] = 8'b00000000;
	mem[1608] = 8'b00000000;
	mem[1609] = 8'b00000000;
	mem[1610] = 8'b00000000;
	mem[1611] = 8'b00000000;
	mem[1612] = 8'b00000000;
	mem[1613] = 8'b00000000;
	mem[1614] = 8'b00000000;
	mem[1615] = 8'b00000000;
	mem[1616] = 8'b00000000;
	mem[1617] = 8'b00000000;
	mem[1618] = 8'b00000000;
	mem[1619] = 8'b00000000;
	mem[1620] = 8'b00000000;
	mem[1621] = 8'b00000000;
	mem[1622] = 8'b00000000;
	mem[1623] = 8'b00000000;
	mem[1624] = 8'b00000000;
	mem[1625] = 8'b00000000;
	mem[1626] = 8'b00000000;
	mem[1627] = 8'b00000000;
	mem[1628] = 8'b00000000;
	mem[1629] = 8'b00000000;
	mem[1630] = 8'b00000000;
	mem[1631] = 8'b00000000;
	mem[1632] = 8'b00000000;
	mem[1633] = 8'b00000000;
	mem[1634] = 8'b00000000;
	mem[1635] = 8'b00000000;
	mem[1636] = 8'b00000000;
	mem[1637] = 8'b00000000;
	mem[1638] = 8'b00000000;
	mem[1639] = 8'b00000000;
	mem[1640] = 8'b00000000;
	mem[1641] = 8'b00000000;
	mem[1642] = 8'b00000000;
	mem[1643] = 8'b00000000;
	mem[1644] = 8'b00000000;
	mem[1645] = 8'b00000000;
	mem[1646] = 8'b00000000;
	mem[1647] = 8'b00000000;
	mem[1648] = 8'b00000000;
	mem[1649] = 8'b00000000;
	mem[1650] = 8'b00000000;
	mem[1651] = 8'b00000000;
	mem[1652] = 8'b00000000;
	mem[1653] = 8'b00000000;
	mem[1654] = 8'b00000000;
	mem[1655] = 8'b00000000;
	mem[1656] = 8'b00000000;
	mem[1657] = 8'b00000000;
	mem[1658] = 8'b00000000;
	mem[1659] = 8'b00000000;
	mem[1660] = 8'b00000000;
	mem[1661] = 8'b00000000;
	mem[1662] = 8'b00000000;
	mem[1663] = 8'b00000000;
	mem[1664] = 8'b00000000;
	mem[1665] = 8'b00000000;
	mem[1666] = 8'b00000000;
	mem[1667] = 8'b00000000;
	mem[1668] = 8'b00000000;
	mem[1669] = 8'b00000000;
	mem[1670] = 8'b00000000;
	mem[1671] = 8'b00000000;
	mem[1672] = 8'b00000000;
	mem[1673] = 8'b00000000;
	mem[1674] = 8'b00000000;
	mem[1675] = 8'b00000000;
	mem[1676] = 8'b00000000;
	mem[1677] = 8'b00000000;
	mem[1678] = 8'b00000000;
	mem[1679] = 8'b00000000;
	mem[1680] = 8'b00000000;
	mem[1681] = 8'b00000000;
	mem[1682] = 8'b00000000;
	mem[1683] = 8'b00000000;
	mem[1684] = 8'b00000000;
	mem[1685] = 8'b00000000;
	mem[1686] = 8'b00000000;
	mem[1687] = 8'b00000000;
	mem[1688] = 8'b00000000;
	mem[1689] = 8'b00000000;
	mem[1690] = 8'b00000000;
	mem[1691] = 8'b00000000;
	mem[1692] = 8'b00000000;
	mem[1693] = 8'b00000000;
	mem[1694] = 8'b00000000;
	mem[1695] = 8'b00000000;
	mem[1696] = 8'b00000000;
	mem[1697] = 8'b00000000;
	mem[1698] = 8'b00000000;
	mem[1699] = 8'b00000000;
	mem[1700] = 8'b00000000;
	mem[1701] = 8'b00000000;
	mem[1702] = 8'b00000000;
	mem[1703] = 8'b00000000;
	mem[1704] = 8'b00000000;
	mem[1705] = 8'b00000000;
	mem[1706] = 8'b00000000;
	mem[1707] = 8'b00000000;
	mem[1708] = 8'b00000000;
	mem[1709] = 8'b00000000;
	mem[1710] = 8'b00000000;
	mem[1711] = 8'b00000000;
	mem[1712] = 8'b00000000;
	mem[1713] = 8'b00000000;
	mem[1714] = 8'b00000000;
	mem[1715] = 8'b00000000;
	mem[1716] = 8'b00000000;
	mem[1717] = 8'b00000000;
	mem[1718] = 8'b00000000;
	mem[1719] = 8'b00000000;
	mem[1720] = 8'b00000000;
	mem[1721] = 8'b00000000;
	mem[1722] = 8'b00000000;
	mem[1723] = 8'b00000000;
	mem[1724] = 8'b00000000;
	mem[1725] = 8'b00000000;
	mem[1726] = 8'b00000000;
	mem[1727] = 8'b00000000;
	mem[1728] = 8'b00000000;
	mem[1729] = 8'b00000000;
	mem[1730] = 8'b00000000;
	mem[1731] = 8'b00000000;
	mem[1732] = 8'b00000000;
	mem[1733] = 8'b00000000;
	mem[1734] = 8'b00000000;
	mem[1735] = 8'b00000000;
	mem[1736] = 8'b00000000;
	mem[1737] = 8'b00000000;
	mem[1738] = 8'b00000000;
	mem[1739] = 8'b00000000;
	mem[1740] = 8'b00000000;
	mem[1741] = 8'b00000000;
	mem[1742] = 8'b00000000;
	mem[1743] = 8'b00000000;
	mem[1744] = 8'b00000000;
	mem[1745] = 8'b00000000;
	mem[1746] = 8'b00000000;
	mem[1747] = 8'b00000000;
	mem[1748] = 8'b00000000;
	mem[1749] = 8'b00000000;
	mem[1750] = 8'b00000000;
	mem[1751] = 8'b00000000;
	mem[1752] = 8'b00000000;
	mem[1753] = 8'b00000000;
	mem[1754] = 8'b00000000;
	mem[1755] = 8'b00000000;
	mem[1756] = 8'b00000000;
	mem[1757] = 8'b00000000;
	mem[1758] = 8'b00000000;
	mem[1759] = 8'b00000000;
	mem[1760] = 8'b00000000;
	mem[1761] = 8'b00000000;
	mem[1762] = 8'b00000000;
	mem[1763] = 8'b00000000;
	mem[1764] = 8'b00000000;
	mem[1765] = 8'b00000000;
	mem[1766] = 8'b00000000;
	mem[1767] = 8'b00000000;
	mem[1768] = 8'b00000000;
	mem[1769] = 8'b00000000;
	mem[1770] = 8'b00000000;
	mem[1771] = 8'b00000000;
	mem[1772] = 8'b00000000;
	mem[1773] = 8'b00000000;
	mem[1774] = 8'b00000000;
	mem[1775] = 8'b00000000;
	mem[1776] = 8'b00000000;
	mem[1777] = 8'b00000000;
	mem[1778] = 8'b00000000;
	mem[1779] = 8'b00000000;
	mem[1780] = 8'b00000000;
	mem[1781] = 8'b00000000;
	mem[1782] = 8'b00000000;
	mem[1783] = 8'b00000000;
	mem[1784] = 8'b00000000;
	mem[1785] = 8'b00000000;
	mem[1786] = 8'b00000000;
	mem[1787] = 8'b00000000;
	mem[1788] = 8'b00000000;
	mem[1789] = 8'b00000000;
	mem[1790] = 8'b00000000;
	mem[1791] = 8'b00000000;
	mem[1792] = 8'b00000000;
	mem[1793] = 8'b00000000;
	mem[1794] = 8'b00000000;
	mem[1795] = 8'b00000000;
	mem[1796] = 8'b00000000;
	mem[1797] = 8'b00000000;
	mem[1798] = 8'b00000000;
	mem[1799] = 8'b00000000;
	mem[1800] = 8'b00000000;
	mem[1801] = 8'b00000000;
	mem[1802] = 8'b00000000;
	mem[1803] = 8'b00000000;
	mem[1804] = 8'b00000000;
	mem[1805] = 8'b00000000;
	mem[1806] = 8'b00000000;
	mem[1807] = 8'b00000000;
	mem[1808] = 8'b00000000;
	mem[1809] = 8'b00000000;
	mem[1810] = 8'b00000000;
	mem[1811] = 8'b00000000;
	mem[1812] = 8'b00000000;
	mem[1813] = 8'b00000000;
	mem[1814] = 8'b00000000;
	mem[1815] = 8'b00000000;
	mem[1816] = 8'b00000000;
	mem[1817] = 8'b00000000;
	mem[1818] = 8'b00000000;
	mem[1819] = 8'b00000000;
	mem[1820] = 8'b00000000;
	mem[1821] = 8'b00000000;
	mem[1822] = 8'b00000000;
	mem[1823] = 8'b00000000;
	mem[1824] = 8'b00000000;
	mem[1825] = 8'b00000000;
	mem[1826] = 8'b00000000;
	mem[1827] = 8'b00000000;
	mem[1828] = 8'b00000000;
	mem[1829] = 8'b00000000;
	mem[1830] = 8'b00000000;
	mem[1831] = 8'b00000000;
	mem[1832] = 8'b00000000;
	mem[1833] = 8'b00000000;
	mem[1834] = 8'b00000000;
	mem[1835] = 8'b00000000;
	mem[1836] = 8'b00000000;
	mem[1837] = 8'b00000000;
	mem[1838] = 8'b00000000;
	mem[1839] = 8'b00000000;
	mem[1840] = 8'b00000000;
	mem[1841] = 8'b00000000;
	mem[1842] = 8'b00000000;
	mem[1843] = 8'b00000000;
	mem[1844] = 8'b00000000;
	mem[1845] = 8'b00000000;
	mem[1846] = 8'b00000000;
	mem[1847] = 8'b00000000;
	mem[1848] = 8'b00000000;
	mem[1849] = 8'b00000000;
	mem[1850] = 8'b00000000;
	mem[1851] = 8'b00000000;
	mem[1852] = 8'b00000000;
	mem[1853] = 8'b00000000;
	mem[1854] = 8'b00000000;
	mem[1855] = 8'b00000000;
	mem[1856] = 8'b00000000;
	mem[1857] = 8'b00000000;
	mem[1858] = 8'b00000000;
	mem[1859] = 8'b00000000;
	mem[1860] = 8'b00000000;
	mem[1861] = 8'b00000000;
	mem[1862] = 8'b00000000;
	mem[1863] = 8'b00000000;
	mem[1864] = 8'b00000000;
	mem[1865] = 8'b00000000;
	mem[1866] = 8'b00000000;
	mem[1867] = 8'b00000000;
	mem[1868] = 8'b00000000;
	mem[1869] = 8'b00000000;
	mem[1870] = 8'b00000000;
	mem[1871] = 8'b00000000;
	mem[1872] = 8'b00000000;
	mem[1873] = 8'b00000000;
	mem[1874] = 8'b00000000;
	mem[1875] = 8'b00000000;
	mem[1876] = 8'b00000000;
	mem[1877] = 8'b00000000;
	mem[1878] = 8'b00000000;
	mem[1879] = 8'b00000000;
	mem[1880] = 8'b00000000;
	mem[1881] = 8'b00000000;
	mem[1882] = 8'b00000000;
	mem[1883] = 8'b00000000;
	mem[1884] = 8'b00000000;
	mem[1885] = 8'b00000000;
	mem[1886] = 8'b00000000;
	mem[1887] = 8'b00000000;
	mem[1888] = 8'b00000000;
	mem[1889] = 8'b00000000;
	mem[1890] = 8'b00000000;
	mem[1891] = 8'b00000000;
	mem[1892] = 8'b00000000;
	mem[1893] = 8'b00000000;
	mem[1894] = 8'b00000000;
	mem[1895] = 8'b00000000;
	mem[1896] = 8'b00000000;
	mem[1897] = 8'b00000000;
	mem[1898] = 8'b00000000;
	mem[1899] = 8'b00000000;
	mem[1900] = 8'b00000000;
	mem[1901] = 8'b00000000;
	mem[1902] = 8'b00000000;
	mem[1903] = 8'b00000000;
	mem[1904] = 8'b00000000;
	mem[1905] = 8'b00000000;
	mem[1906] = 8'b00000000;
	mem[1907] = 8'b00000000;
	mem[1908] = 8'b00000000;
	mem[1909] = 8'b00000000;
	mem[1910] = 8'b00000000;
	mem[1911] = 8'b00000000;
	mem[1912] = 8'b00000000;
	mem[1913] = 8'b00000000;
	mem[1914] = 8'b00000000;
	mem[1915] = 8'b00000000;
	mem[1916] = 8'b00000000;
	mem[1917] = 8'b00000000;
	mem[1918] = 8'b00000000;
	mem[1919] = 8'b00000000;
	mem[1920] = 8'b00000000;
	mem[1921] = 8'b00000000;
	mem[1922] = 8'b00000000;
	mem[1923] = 8'b00000000;
	mem[1924] = 8'b00000000;
	mem[1925] = 8'b00000000;
	mem[1926] = 8'b00000000;
	mem[1927] = 8'b00000000;
	mem[1928] = 8'b00000000;
	mem[1929] = 8'b00000000;
	mem[1930] = 8'b00000000;
	mem[1931] = 8'b00000000;
	mem[1932] = 8'b00000000;
	mem[1933] = 8'b00000000;
	mem[1934] = 8'b00000000;
	mem[1935] = 8'b00000000;
	mem[1936] = 8'b00000000;
	mem[1937] = 8'b00000000;
	mem[1938] = 8'b00000000;
	mem[1939] = 8'b00000000;
	mem[1940] = 8'b00000000;
	mem[1941] = 8'b00000000;
	mem[1942] = 8'b00000000;
	mem[1943] = 8'b00000000;
	mem[1944] = 8'b00000000;
	mem[1945] = 8'b00000000;
	mem[1946] = 8'b00000000;
	mem[1947] = 8'b00000000;
	mem[1948] = 8'b00000000;
	mem[1949] = 8'b00000000;
	mem[1950] = 8'b00000000;
	mem[1951] = 8'b00000000;
	mem[1952] = 8'b00000000;
	mem[1953] = 8'b00000000;
	mem[1954] = 8'b00000000;
	mem[1955] = 8'b00000000;
	mem[1956] = 8'b00000000;
	mem[1957] = 8'b00000000;
	mem[1958] = 8'b00000000;
	mem[1959] = 8'b00000000;
	mem[1960] = 8'b00000000;
	mem[1961] = 8'b00000000;
	mem[1962] = 8'b00000000;
	mem[1963] = 8'b00000000;
	mem[1964] = 8'b00000000;
	mem[1965] = 8'b00000000;
	mem[1966] = 8'b00000000;
	mem[1967] = 8'b00000000;
	mem[1968] = 8'b00000000;
	mem[1969] = 8'b00000000;
	mem[1970] = 8'b00000000;
	mem[1971] = 8'b00000000;
	mem[1972] = 8'b00000000;
	mem[1973] = 8'b00000000;
	mem[1974] = 8'b00000000;
	mem[1975] = 8'b00000000;
	mem[1976] = 8'b00000000;
	mem[1977] = 8'b00000000;
	mem[1978] = 8'b00000000;
	mem[1979] = 8'b00000000;
	mem[1980] = 8'b00000000;
	mem[1981] = 8'b00000000;
	mem[1982] = 8'b00000000;
	mem[1983] = 8'b00000000;
	mem[1984] = 8'b00000000;
	mem[1985] = 8'b00000000;
	mem[1986] = 8'b00000000;
	mem[1987] = 8'b00000000;
	mem[1988] = 8'b00000000;
	mem[1989] = 8'b00000000;
	mem[1990] = 8'b00000000;
	mem[1991] = 8'b00000000;
	mem[1992] = 8'b00000000;
	mem[1993] = 8'b00000000;
	mem[1994] = 8'b00000000;
	mem[1995] = 8'b00000000;
	mem[1996] = 8'b00000000;
	mem[1997] = 8'b00000000;
	mem[1998] = 8'b00000000;
	mem[1999] = 8'b00000000;
	mem[2000] = 8'b00000000;
	mem[2001] = 8'b00000000;
	mem[2002] = 8'b00000000;
	mem[2003] = 8'b00000000;
	mem[2004] = 8'b00000000;
	mem[2005] = 8'b00000000;
	mem[2006] = 8'b00000000;
	mem[2007] = 8'b00000000;
	mem[2008] = 8'b00000000;
	mem[2009] = 8'b00000000;
	mem[2010] = 8'b00000000;
	mem[2011] = 8'b00000000;
	mem[2012] = 8'b00000000;
	mem[2013] = 8'b00000000;
	mem[2014] = 8'b00000000;
	mem[2015] = 8'b00000000;
	mem[2016] = 8'b00000000;
	mem[2017] = 8'b00000000;
	mem[2018] = 8'b00000000;
	mem[2019] = 8'b00000000;
	mem[2020] = 8'b00000000;
	mem[2021] = 8'b00000000;
	mem[2022] = 8'b00000000;
	mem[2023] = 8'b00000000;
	mem[2024] = 8'b00000000;
	mem[2025] = 8'b00000000;
	mem[2026] = 8'b00000000;
	mem[2027] = 8'b00000000;
	mem[2028] = 8'b00000000;
	mem[2029] = 8'b00000000;
	mem[2030] = 8'b00000000;
	mem[2031] = 8'b00000000;
	mem[2032] = 8'b00000000;
	mem[2033] = 8'b00000000;
	mem[2034] = 8'b00000000;
	mem[2035] = 8'b00000000;
	mem[2036] = 8'b00000000;
	mem[2037] = 8'b00000000;
	mem[2038] = 8'b00000000;
	mem[2039] = 8'b00000000;
	mem[2040] = 8'b00000000;
	mem[2041] = 8'b00000000;
	mem[2042] = 8'b00000000;
	mem[2043] = 8'b00000000;
	mem[2044] = 8'b00000000;
	mem[2045] = 8'b00000000;
	mem[2046] = 8'b00000000;
	mem[2047] = 8'b00000000;
end
endmodule
