module char_rom_r(
	input clock,
	input [8:0] address,
	output reg [7:0] data_out
);

reg [7:0] mem [0:511];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 8'b00001111;
	mem[1] = 8'b00001111;
	mem[2] = 8'b00001111;
	mem[3] = 8'b00001101;
	mem[4] = 8'b00001011;
	mem[5] = 8'b00001011;
	mem[6] = 8'b00001101;
	mem[7] = 8'b00001101;
	mem[8] = 8'b00001101;
	mem[9] = 8'b00001011;
	mem[10] = 8'b00001111;
	mem[11] = 8'b00001111;
	mem[12] = 8'b00001111;
	mem[13] = 8'b00001100;
	mem[14] = 8'b00001100;
	mem[15] = 8'b00001011;
	mem[16] = 8'b00001111;
	mem[17] = 8'b00001111;
	mem[18] = 8'b00001111;
	mem[19] = 8'b00001011;
	mem[20] = 8'b00001011;
	mem[21] = 8'b00001100;
	mem[22] = 8'b00001111;
	mem[23] = 8'b00001111;
	mem[24] = 8'b00001111;
	mem[25] = 8'b00001111;
	mem[26] = 8'b00001110;
	mem[27] = 8'b00001011;
	mem[28] = 8'b00001011;
	mem[29] = 8'b00001100;
	mem[30] = 8'b00001111;
	mem[31] = 8'b00001111;
	mem[32] = 8'b00001100;
	mem[33] = 8'b00001100;
	mem[34] = 8'b00001100;
	mem[35] = 8'b00001101;
	mem[36] = 8'b00001111;
	mem[37] = 8'b00001111;
	mem[38] = 8'b00001111;
	mem[39] = 8'b00001101;
	mem[40] = 8'b00001110;
	mem[41] = 8'b00001111;
	mem[42] = 8'b00001111;
	mem[43] = 8'b00001111;
	mem[44] = 8'b00001111;
	mem[45] = 8'b00001111;
	mem[46] = 8'b00001111;
	mem[47] = 8'b00001111;
	mem[48] = 8'b00001111;
	mem[49] = 8'b00001111;
	mem[50] = 8'b00001111;
	mem[51] = 8'b00001111;
	mem[52] = 8'b00001111;
	mem[53] = 8'b00001111;
	mem[54] = 8'b00001111;
	mem[55] = 8'b00001111;
	mem[56] = 8'b00001111;
	mem[57] = 8'b00001111;
	mem[58] = 8'b00001111;
	mem[59] = 8'b00001111;
	mem[60] = 8'b00001111;
	mem[61] = 8'b00001111;
	mem[62] = 8'b00001111;
	mem[63] = 8'b00001111;
	mem[64] = 8'b00001111;
	mem[65] = 8'b00001110;
	mem[66] = 8'b00001011;
	mem[67] = 8'b00001111;
	mem[68] = 8'b00001111;
	mem[69] = 8'b00001111;
	mem[70] = 8'b00001101;
	mem[71] = 8'b00001100;
	mem[72] = 8'b00001100;
	mem[73] = 8'b00001011;
	mem[74] = 8'b00001111;
	mem[75] = 8'b00001111;
	mem[76] = 8'b00001011;
	mem[77] = 8'b00001111;
	mem[78] = 8'b00001111;
	mem[79] = 8'b00001011;
	mem[80] = 8'b00001111;
	mem[81] = 8'b00001111;
	mem[82] = 8'b00001011;
	mem[83] = 8'b00001111;
	mem[84] = 8'b00001111;
	mem[85] = 8'b00001101;
	mem[86] = 8'b00001111;
	mem[87] = 8'b00001111;
	mem[88] = 8'b00001111;
	mem[89] = 8'b00001101;
	mem[90] = 8'b00001101;
	mem[91] = 8'b00001111;
	mem[92] = 8'b00001111;
	mem[93] = 8'b00001011;
	mem[94] = 8'b00001111;
	mem[95] = 8'b00001111;
	mem[96] = 8'b00001101;
	mem[97] = 8'b00001111;
	mem[98] = 8'b00001110;
	mem[99] = 8'b00001111;
	mem[100] = 8'b00001101;
	mem[101] = 8'b00001110;
	mem[102] = 8'b00001110;
	mem[103] = 8'b00001111;
	mem[104] = 8'b00001110;
	mem[105] = 8'b00001100;
	mem[106] = 8'b00001101;
	mem[107] = 8'b00001100;
	mem[108] = 8'b00001110;
	mem[109] = 8'b00001011;
	mem[110] = 8'b00001110;
	mem[111] = 8'b00001111;
	mem[112] = 8'b00001011;
	mem[113] = 8'b00001110;
	mem[114] = 8'b00001011;
	mem[115] = 8'b00001011;
	mem[116] = 8'b00001011;
	mem[117] = 8'b00001011;
	mem[118] = 8'b00001011;
	mem[119] = 8'b00001011;
	mem[120] = 8'b00001100;
	mem[121] = 8'b00001111;
	mem[122] = 8'b00001011;
	mem[123] = 8'b00001011;
	mem[124] = 8'b00001100;
	mem[125] = 8'b00001101;
	mem[126] = 8'b00001011;
	mem[127] = 8'b00001100;
	mem[128] = 8'b00001101;
	mem[129] = 8'b00001101;
	mem[130] = 8'b00001111;
	mem[131] = 8'b00001111;
	mem[132] = 8'b00001011;
	mem[133] = 8'b00001101;
	mem[134] = 8'b00001111;
	mem[135] = 8'b00001111;
	mem[136] = 8'b00001111;
	mem[137] = 8'b00001111;
	mem[138] = 8'b00001111;
	mem[139] = 8'b00001111;
	mem[140] = 8'b00001101;
	mem[141] = 8'b00001111;
	mem[142] = 8'b00001110;
	mem[143] = 8'b00001011;
	mem[144] = 8'b00001011;
	mem[145] = 8'b00001011;
	mem[146] = 8'b00001101;
	mem[147] = 8'b00001111;
	mem[148] = 8'b00001100;
	mem[149] = 8'b00001111;
	mem[150] = 8'b00001111;
	mem[151] = 8'b00001111;
	mem[152] = 8'b00001101;
	mem[153] = 8'b00001101;
	mem[154] = 8'b00001111;
	mem[155] = 8'b00001100;
	mem[156] = 8'b00001111;
	mem[157] = 8'b00001011;
	mem[158] = 8'b00001111;
	mem[159] = 8'b00001100;
	mem[160] = 8'b00001111;
	mem[161] = 8'b00001100;
	mem[162] = 8'b00001101;
	mem[163] = 8'b00001100;
	mem[164] = 8'b00001111;
	mem[165] = 8'b00001101;
	mem[166] = 8'b00001011;
	mem[167] = 8'b00001111;
	mem[168] = 8'b00001100;
	mem[169] = 8'b00001110;
	mem[170] = 8'b00001111;
	mem[171] = 8'b00001110;
	mem[172] = 8'b00001110;
	mem[173] = 8'b00001111;
	mem[174] = 8'b00001111;
	mem[175] = 8'b00001100;
	mem[176] = 8'b00001111;
	mem[177] = 8'b00001110;
	mem[178] = 8'b00001101;
	mem[179] = 8'b00001110;
	mem[180] = 8'b00001011;
	mem[181] = 8'b00001101;
	mem[182] = 8'b00001100;
	mem[183] = 8'b00001011;
	mem[184] = 8'b00001110;
	mem[185] = 8'b00001101;
	mem[186] = 8'b00001110;
	mem[187] = 8'b00001011;
	mem[188] = 8'b00001101;
	mem[189] = 8'b00001011;
	mem[190] = 8'b00001011;
	mem[191] = 8'b00001110;
	mem[192] = 8'b00001100;
	mem[193] = 8'b00001111;
	mem[194] = 8'b00001111;
	mem[195] = 8'b00001011;
	mem[196] = 8'b00001111;
	mem[197] = 8'b00001111;
	mem[198] = 8'b00001111;
	mem[199] = 8'b00001111;
	mem[200] = 8'b00001111;
	mem[201] = 8'b00001111;
	mem[202] = 8'b00001111;
	mem[203] = 8'b00001011;
	mem[204] = 8'b00001111;
	mem[205] = 8'b00001111;
	mem[206] = 8'b00001111;
	mem[207] = 8'b00001111;
	mem[208] = 8'b00001111;
	mem[209] = 8'b00001111;
	mem[210] = 8'b00001111;
	mem[211] = 8'b00001111;
	mem[212] = 8'b00001100;
	mem[213] = 8'b00001111;
	mem[214] = 8'b00001111;
	mem[215] = 8'b00001100;
	mem[216] = 8'b00001110;
	mem[217] = 8'b00001111;
	mem[218] = 8'b00001100;
	mem[219] = 8'b00001011;
	mem[220] = 8'b00001111;
	mem[221] = 8'b00001101;
	mem[222] = 8'b00001111;
	mem[223] = 8'b00001100;
	mem[224] = 8'b00001111;
	mem[225] = 8'b00001111;
	mem[226] = 8'b00001111;
	mem[227] = 8'b00001110;
	mem[228] = 8'b00001011;
	mem[229] = 8'b00001111;
	mem[230] = 8'b00001101;
	mem[231] = 8'b00001100;
	mem[232] = 8'b00001111;
	mem[233] = 8'b00001011;
	mem[234] = 8'b00001100;
	mem[235] = 8'b00001101;
	mem[236] = 8'b00001011;
	mem[237] = 8'b00001111;
	mem[238] = 8'b00001101;
	mem[239] = 8'b00001110;
	mem[240] = 8'b00001100;
	mem[241] = 8'b00001100;
	mem[242] = 8'b00001110;
	mem[243] = 8'b00001011;
	mem[244] = 8'b00001110;
	mem[245] = 8'b00001101;
	mem[246] = 8'b00001011;
	mem[247] = 8'b00001101;
	mem[248] = 8'b00001101;
	mem[249] = 8'b00001011;
	mem[250] = 8'b00001101;
	mem[251] = 8'b00001100;
	mem[252] = 8'b00001111;
	mem[253] = 8'b00001110;
	mem[254] = 8'b00001110;
	mem[255] = 8'b00001011;
	mem[256] = 8'b00001101;
	mem[257] = 8'b00001111;
	mem[258] = 8'b00001111;
	mem[259] = 8'b00001011;
	mem[260] = 8'b00001111;
	mem[261] = 8'b00001111;
	mem[262] = 8'b00001111;
	mem[263] = 8'b00001100;
	mem[264] = 8'b00001011;
	mem[265] = 8'b00001111;
	mem[266] = 8'b00001111;
	mem[267] = 8'b00001101;
	mem[268] = 8'b00001111;
	mem[269] = 8'b00001101;
	mem[270] = 8'b00001110;
	mem[271] = 8'b00001110;
	mem[272] = 8'b00001110;
	mem[273] = 8'b00001100;
	mem[274] = 8'b00001111;
	mem[275] = 8'b00001101;
	mem[276] = 8'b00001111;
	mem[277] = 8'b00001111;
	mem[278] = 8'b00001100;
	mem[279] = 8'b00001110;
	mem[280] = 8'b00001111;
	mem[281] = 8'b00001111;
	mem[282] = 8'b00001111;
	mem[283] = 8'b00001111;
	mem[284] = 8'b00001111;
	mem[285] = 8'b00001110;
	mem[286] = 8'b00001101;
	mem[287] = 8'b00001111;
	mem[288] = 8'b00001100;
	mem[289] = 8'b00001110;
	mem[290] = 8'b00001111;
	mem[291] = 8'b00001100;
	mem[292] = 8'b00001111;
	mem[293] = 8'b00001100;
	mem[294] = 8'b00001111;
	mem[295] = 8'b00001011;
	mem[296] = 8'b00001111;
	mem[297] = 8'b00001111;
	mem[298] = 8'b00001100;
	mem[299] = 8'b00001111;
	mem[300] = 8'b00001100;
	mem[301] = 8'b00001110;
	mem[302] = 8'b00001110;
	mem[303] = 8'b00001101;
	mem[304] = 8'b00001100;
	mem[305] = 8'b00001101;
	mem[306] = 8'b00001100;
	mem[307] = 8'b00001101;
	mem[308] = 8'b00001100;
	mem[309] = 8'b00001111;
	mem[310] = 8'b00001011;
	mem[311] = 8'b00001101;
	mem[312] = 8'b00001011;
	mem[313] = 8'b00001100;
	mem[314] = 8'b00001100;
	mem[315] = 8'b00001011;
	mem[316] = 8'b00001011;
	mem[317] = 8'b00001100;
	mem[318] = 8'b00001011;
	mem[319] = 8'b00001100;
	mem[320] = 8'b00001011;
	mem[321] = 8'b00001111;
	mem[322] = 8'b00001111;
	mem[323] = 8'b00001111;
	mem[324] = 8'b00001101;
	mem[325] = 8'b00001101;
	mem[326] = 8'b00001110;
	mem[327] = 8'b00001111;
	mem[328] = 8'b00001111;
	mem[329] = 8'b00001011;
	mem[330] = 8'b00001011;
	mem[331] = 8'b00001111;
	mem[332] = 8'b00001111;
	mem[333] = 8'b00001011;
	mem[334] = 8'b00001111;
	mem[335] = 8'b00001111;
	mem[336] = 8'b00001100;
	mem[337] = 8'b00001111;
	mem[338] = 8'b00001111;
	mem[339] = 8'b00001011;
	mem[340] = 8'b00001111;
	mem[341] = 8'b00001100;
	mem[342] = 8'b00001110;
	mem[343] = 8'b00001111;
	mem[344] = 8'b00001011;
	mem[345] = 8'b00001110;
	mem[346] = 8'b00001110;
	mem[347] = 8'b00001111;
	mem[348] = 8'b00001100;
	mem[349] = 8'b00001111;
	mem[350] = 8'b00001011;
	mem[351] = 8'b00001111;
	mem[352] = 8'b00001011;
	mem[353] = 8'b00001111;
	mem[354] = 8'b00001101;
	mem[355] = 8'b00001110;
	mem[356] = 8'b00001111;
	mem[357] = 8'b00001011;
	mem[358] = 8'b00001110;
	mem[359] = 8'b00001101;
	mem[360] = 8'b00001100;
	mem[361] = 8'b00001100;
	mem[362] = 8'b00001011;
	mem[363] = 8'b00001100;
	mem[364] = 8'b00001100;
	mem[365] = 8'b00001011;
	mem[366] = 8'b00001011;
	mem[367] = 8'b00001100;
	mem[368] = 8'b00001100;
	mem[369] = 8'b00001011;
	mem[370] = 8'b00001011;
	mem[371] = 8'b00001100;
	mem[372] = 8'b00001100;
	mem[373] = 8'b00001011;
	mem[374] = 8'b00001011;
	mem[375] = 8'b00001100;
	mem[376] = 8'b00001101;
	mem[377] = 8'b00001011;
	mem[378] = 8'b00001100;
	mem[379] = 8'b00001100;
	mem[380] = 8'b00001110;
	mem[381] = 8'b00001110;
	mem[382] = 8'b00001101;
	mem[383] = 8'b00001110;
	mem[384] = 8'b00001111;
	mem[385] = 8'b00001101;
	mem[386] = 8'b00001011;
	mem[387] = 8'b00001100;
	mem[388] = 8'b00001100;
	mem[389] = 8'b00001100;
	mem[390] = 8'b00001100;
	mem[391] = 8'b00001011;
	mem[392] = 8'b00001100;
	mem[393] = 8'b00001111;
	mem[394] = 8'b00001011;
	mem[395] = 8'b00001100;
	mem[396] = 8'b00001101;
	mem[397] = 8'b00001111;
	mem[398] = 8'b00001111;
	mem[399] = 8'b00001111;
	mem[400] = 8'b00001100;
	mem[401] = 8'b00001011;
	mem[402] = 8'b00001011;
	mem[403] = 8'b00001111;
	mem[404] = 8'b00001111;
	mem[405] = 8'b00001111;
	mem[406] = 8'b00001011;
	mem[407] = 8'b00001100;
	mem[408] = 8'b00001111;
	mem[409] = 8'b00001111;
	mem[410] = 8'b00001111;
	mem[411] = 8'b00001111;
	mem[412] = 8'b00001101;
	mem[413] = 8'b00001110;
	mem[414] = 8'b00001111;
	mem[415] = 8'b00001111;
	mem[416] = 8'b00001111;
	mem[417] = 8'b00001111;
	mem[418] = 8'b00001110;
	mem[419] = 8'b00001111;
	mem[420] = 8'b00001111;
	mem[421] = 8'b00001111;
	mem[422] = 8'b00001111;
	mem[423] = 8'b00001111;
	mem[424] = 8'b00001111;
	mem[425] = 8'b00001111;
	mem[426] = 8'b00001111;
	mem[427] = 8'b00001111;
	mem[428] = 8'b00001111;
	mem[429] = 8'b00001111;
	mem[430] = 8'b00001111;
	mem[431] = 8'b00001111;
	mem[432] = 8'b00001111;
	mem[433] = 8'b00001111;
	mem[434] = 8'b00001111;
	mem[435] = 8'b00001111;
	mem[436] = 8'b00001111;
	mem[437] = 8'b00001111;
	mem[438] = 8'b00001111;
	mem[439] = 8'b00001111;
	mem[440] = 8'b00001111;
	mem[441] = 8'b00001111;
	mem[442] = 8'b00001111;
	mem[443] = 8'b00001111;
	mem[444] = 8'b00001111;
	mem[445] = 8'b00001111;
	mem[446] = 8'b00001111;
	mem[447] = 8'b00001111;
	mem[448] = 8'b00000000;
	mem[449] = 8'b00000000;
	mem[450] = 8'b00000000;
	mem[451] = 8'b00000000;
	mem[452] = 8'b00000000;
	mem[453] = 8'b00000000;
	mem[454] = 8'b00000000;
	mem[455] = 8'b00000000;
	mem[456] = 8'b00000000;
	mem[457] = 8'b00000000;
	mem[458] = 8'b00000000;
	mem[459] = 8'b00000000;
	mem[460] = 8'b00000000;
	mem[461] = 8'b00000000;
	mem[462] = 8'b00000000;
	mem[463] = 8'b00000000;
	mem[464] = 8'b00000000;
	mem[465] = 8'b00000000;
	mem[466] = 8'b00000000;
	mem[467] = 8'b00000000;
	mem[468] = 8'b00000000;
	mem[469] = 8'b00000000;
	mem[470] = 8'b00000000;
	mem[471] = 8'b00000000;
	mem[472] = 8'b00000000;
	mem[473] = 8'b00000000;
	mem[474] = 8'b00000000;
	mem[475] = 8'b00000000;
	mem[476] = 8'b00000000;
	mem[477] = 8'b00000000;
	mem[478] = 8'b00000000;
	mem[479] = 8'b00000000;
	mem[480] = 8'b00000000;
	mem[481] = 8'b00000000;
	mem[482] = 8'b00000000;
	mem[483] = 8'b00000000;
	mem[484] = 8'b00000000;
	mem[485] = 8'b00000000;
	mem[486] = 8'b00000000;
	mem[487] = 8'b00000000;
	mem[488] = 8'b00000000;
	mem[489] = 8'b00000000;
	mem[490] = 8'b00000000;
	mem[491] = 8'b00000000;
	mem[492] = 8'b00000000;
	mem[493] = 8'b00000000;
	mem[494] = 8'b00000000;
	mem[495] = 8'b00000000;
	mem[496] = 8'b00000000;
	mem[497] = 8'b00000000;
	mem[498] = 8'b00000000;
	mem[499] = 8'b00000000;
	mem[500] = 8'b00000000;
	mem[501] = 8'b00000000;
	mem[502] = 8'b00000000;
	mem[503] = 8'b00000000;
	mem[504] = 8'b00000000;
	mem[505] = 8'b00000000;
	mem[506] = 8'b00000000;
	mem[507] = 8'b00000000;
	mem[508] = 8'b00000000;
	mem[509] = 8'b00000000;
	mem[510] = 8'b00000000;
	mem[511] = 8'b00000000;
end
endmodule
